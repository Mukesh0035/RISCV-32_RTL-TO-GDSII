magic
tech sky130A
magscale 1 2
timestamp 1753979594
<< checkpaint >>
rect -3932 -3932 15122 17266
<< viali >>
rect 2237 10761 2271 10795
rect 2789 10761 2823 10795
rect 4169 10761 4203 10795
rect 6469 10761 6503 10795
rect 7297 10761 7331 10795
rect 9321 10761 9355 10795
rect 1777 10625 1811 10659
rect 2329 10625 2363 10659
rect 3065 10625 3099 10659
rect 3433 10625 3467 10659
rect 4077 10625 4111 10659
rect 6745 10625 6779 10659
rect 7573 10625 7607 10659
rect 9045 10625 9079 10659
rect 8493 10557 8527 10591
rect 1501 10421 1535 10455
rect 3249 10421 3283 10455
rect 7941 10421 7975 10455
rect 3341 10217 3375 10251
rect 3801 10217 3835 10251
rect 9597 10217 9631 10251
rect 3065 10149 3099 10183
rect 4353 10081 4387 10115
rect 7389 10081 7423 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 4905 10013 4939 10047
rect 5457 10013 5491 10047
rect 7021 10013 7055 10047
rect 7113 10013 7147 10047
rect 9137 10013 9171 10047
rect 1952 9945 1986 9979
rect 3249 9945 3283 9979
rect 4997 9945 5031 9979
rect 5181 9945 5215 9979
rect 5724 9945 5758 9979
rect 7656 9945 7690 9979
rect 9321 9945 9355 9979
rect 1593 9877 1627 9911
rect 4721 9877 4755 9911
rect 5365 9877 5399 9911
rect 6837 9877 6871 9911
rect 7297 9877 7331 9911
rect 8769 9877 8803 9911
rect 8953 9877 8987 9911
rect 2237 9673 2271 9707
rect 3617 9673 3651 9707
rect 5825 9673 5859 9707
rect 1593 9605 1627 9639
rect 6377 9605 6411 9639
rect 7297 9605 7331 9639
rect 8576 9605 8610 9639
rect 1961 9537 1995 9571
rect 2421 9537 2455 9571
rect 3433 9537 3467 9571
rect 4721 9537 4755 9571
rect 5089 9537 5123 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 7481 9537 7515 9571
rect 8125 9537 8159 9571
rect 3065 9469 3099 9503
rect 7021 9469 7055 9503
rect 8309 9469 8343 9503
rect 5089 9401 5123 9435
rect 9689 9401 9723 9435
rect 2513 9333 2547 9367
rect 5365 9333 5399 9367
rect 7113 9333 7147 9367
rect 8033 9333 8067 9367
rect 3341 9129 3375 9163
rect 7573 9129 7607 9163
rect 7941 9129 7975 9163
rect 8217 9129 8251 9163
rect 1593 8993 1627 9027
rect 9689 8993 9723 9027
rect 3617 8925 3651 8959
rect 5825 8925 5859 8959
rect 7849 8925 7883 8959
rect 8125 8925 8159 8959
rect 8401 8925 8435 8959
rect 8493 8925 8527 8959
rect 1869 8857 1903 8891
rect 3525 8857 3559 8891
rect 6101 8857 6135 8891
rect 7757 8857 7791 8891
rect 8677 8789 8711 8823
rect 9045 8789 9079 8823
rect 2329 8585 2363 8619
rect 9229 8585 9263 8619
rect 4721 8517 4755 8551
rect 1593 8449 1627 8483
rect 2421 8449 2455 8483
rect 2605 8449 2639 8483
rect 2697 8449 2731 8483
rect 4813 8449 4847 8483
rect 5080 8449 5114 8483
rect 8861 8449 8895 8483
rect 9505 8449 9539 8483
rect 1685 8381 1719 8415
rect 1961 8381 1995 8415
rect 2973 8381 3007 8415
rect 6193 8313 6227 8347
rect 9045 8313 9079 8347
rect 1501 8041 1535 8075
rect 3341 8041 3375 8075
rect 3893 8041 3927 8075
rect 4997 8041 5031 8075
rect 6193 8041 6227 8075
rect 2053 7905 2087 7939
rect 4077 7905 4111 7939
rect 4721 7905 4755 7939
rect 6929 7905 6963 7939
rect 7021 7905 7055 7939
rect 1777 7837 1811 7871
rect 2145 7837 2179 7871
rect 2973 7837 3007 7871
rect 3433 7837 3467 7871
rect 3985 7837 4019 7871
rect 4813 7837 4847 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 6745 7837 6779 7871
rect 7113 7837 7147 7871
rect 7297 7837 7331 7871
rect 8125 7837 8159 7871
rect 2789 7769 2823 7803
rect 9321 7769 9355 7803
rect 3157 7701 3191 7735
rect 6561 7701 6595 7735
rect 8309 7701 8343 7735
rect 9597 7701 9631 7735
rect 2881 7497 2915 7531
rect 5089 7497 5123 7531
rect 6653 7497 6687 7531
rect 9689 7497 9723 7531
rect 4353 7429 4387 7463
rect 5273 7429 5307 7463
rect 8554 7429 8588 7463
rect 4905 7361 4939 7395
rect 5457 7361 5491 7395
rect 6745 7361 6779 7395
rect 7389 7361 7423 7395
rect 7665 7361 7699 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 4629 7293 4663 7327
rect 4721 7293 4755 7327
rect 4813 7293 4847 7327
rect 6469 7293 6503 7327
rect 7573 7293 7607 7327
rect 4445 7157 4479 7191
rect 7113 7157 7147 7191
rect 7205 7157 7239 7191
rect 8125 7157 8159 7191
rect 2421 6953 2455 6987
rect 7757 6953 7791 6987
rect 8033 6953 8067 6987
rect 8953 6953 8987 6987
rect 2789 6817 2823 6851
rect 3525 6817 3559 6851
rect 6469 6817 6503 6851
rect 6745 6817 6779 6851
rect 7021 6817 7055 6851
rect 8769 6817 8803 6851
rect 9137 6817 9171 6851
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 2145 6749 2179 6783
rect 2697 6749 2731 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 3157 6749 3191 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 4353 6749 4387 6783
rect 4629 6749 4663 6783
rect 7113 6749 7147 6783
rect 7481 6749 7515 6783
rect 7849 6749 7883 6783
rect 9229 6749 9263 6783
rect 1409 6681 1443 6715
rect 1777 6681 1811 6715
rect 2605 6681 2639 6715
rect 3801 6681 3835 6715
rect 4905 6681 4939 6715
rect 8125 6681 8159 6715
rect 9597 6681 9631 6715
rect 2237 6613 2271 6647
rect 2405 6613 2439 6647
rect 4721 6613 4755 6647
rect 3157 6409 3191 6443
rect 4537 6409 4571 6443
rect 6929 6409 6963 6443
rect 7849 6409 7883 6443
rect 9505 6409 9539 6443
rect 1685 6341 1719 6375
rect 3617 6341 3651 6375
rect 3433 6273 3467 6307
rect 3985 6273 4019 6307
rect 4169 6273 4203 6307
rect 4445 6273 4479 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 8381 6273 8415 6307
rect 1409 6205 1443 6239
rect 3249 6205 3283 6239
rect 4813 6205 4847 6239
rect 5457 6205 5491 6239
rect 8125 6205 8159 6239
rect 3893 6069 3927 6103
rect 4261 6069 4295 6103
rect 4997 6069 5031 6103
rect 5273 6069 5307 6103
rect 5733 6069 5767 6103
rect 2237 5865 2271 5899
rect 4261 5865 4295 5899
rect 4997 5865 5031 5899
rect 5181 5865 5215 5899
rect 6653 5865 6687 5899
rect 7297 5729 7331 5763
rect 8953 5729 8987 5763
rect 9505 5729 9539 5763
rect 3361 5661 3395 5695
rect 3617 5661 3651 5695
rect 5917 5661 5951 5695
rect 6009 5661 6043 5695
rect 6285 5661 6319 5695
rect 6377 5661 6411 5695
rect 7021 5661 7055 5695
rect 7481 5661 7515 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 1777 5593 1811 5627
rect 4077 5593 4111 5627
rect 4813 5593 4847 5627
rect 5013 5593 5047 5627
rect 6101 5593 6135 5627
rect 1869 5525 1903 5559
rect 4277 5525 4311 5559
rect 4445 5525 4479 5559
rect 5733 5525 5767 5559
rect 6469 5525 6503 5559
rect 6653 5525 6687 5559
rect 8033 5525 8067 5559
rect 4353 5321 4387 5355
rect 6377 5321 6411 5355
rect 6561 5321 6595 5355
rect 9321 5321 9355 5355
rect 8186 5253 8220 5287
rect 9413 5253 9447 5287
rect 9597 5253 9631 5287
rect 2329 5185 2363 5219
rect 2605 5185 2639 5219
rect 3893 5185 3927 5219
rect 4721 5185 4755 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 5733 5185 5767 5219
rect 6929 5185 6963 5219
rect 7021 5185 7055 5219
rect 7205 5185 7239 5219
rect 7481 5185 7515 5219
rect 7941 5185 7975 5219
rect 1685 5117 1719 5151
rect 5641 5117 5675 5151
rect 6101 5117 6135 5151
rect 7389 5117 7423 5151
rect 7573 5117 7607 5151
rect 7665 5117 7699 5151
rect 7113 5049 7147 5083
rect 2421 4981 2455 5015
rect 3985 4981 4019 5015
rect 4905 4981 4939 5015
rect 5365 4981 5399 5015
rect 6561 4981 6595 5015
rect 7849 4981 7883 5015
rect 1409 4777 1443 4811
rect 7849 4777 7883 4811
rect 9045 4777 9079 4811
rect 4629 4709 4663 4743
rect 5181 4641 5215 4675
rect 7021 4641 7055 4675
rect 7389 4641 7423 4675
rect 2789 4573 2823 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5365 4573 5399 4607
rect 7205 4573 7239 4607
rect 7665 4573 7699 4607
rect 9597 4573 9631 4607
rect 2522 4505 2556 4539
rect 5273 4505 5307 4539
rect 7481 4505 7515 4539
rect 8401 4505 8435 4539
rect 8769 4505 8803 4539
rect 5089 4437 5123 4471
rect 4721 4233 4755 4267
rect 5365 4233 5399 4267
rect 9689 4233 9723 4267
rect 2237 4165 2271 4199
rect 1501 4097 1535 4131
rect 1777 4097 1811 4131
rect 2421 4097 2455 4131
rect 2697 4097 2731 4131
rect 4353 4097 4387 4131
rect 5181 4097 5215 4131
rect 5457 4097 5491 4131
rect 6929 4097 6963 4131
rect 7113 4097 7147 4131
rect 8309 4097 8343 4131
rect 8565 4097 8599 4131
rect 2053 4029 2087 4063
rect 2881 4029 2915 4063
rect 3525 4029 3559 4063
rect 4445 4029 4479 4063
rect 6101 4029 6135 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 1685 3893 1719 3927
rect 1961 3893 1995 3927
rect 2513 3893 2547 3927
rect 4997 3893 5031 3927
rect 5549 3893 5583 3927
rect 7297 3893 7331 3927
rect 4077 3689 4111 3723
rect 7021 3689 7055 3723
rect 3801 3621 3835 3655
rect 5549 3621 5583 3655
rect 2145 3553 2179 3587
rect 2401 3485 2435 3519
rect 3985 3485 4019 3519
rect 4256 3485 4290 3519
rect 4445 3485 4479 3519
rect 4573 3485 4607 3519
rect 4721 3485 4755 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5273 3485 5307 3519
rect 5365 3485 5399 3519
rect 5641 3485 5675 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7757 3485 7791 3519
rect 8953 3485 8987 3519
rect 9505 3485 9539 3519
rect 1777 3417 1811 3451
rect 4353 3417 4387 3451
rect 5886 3417 5920 3451
rect 7665 3417 7699 3451
rect 8401 3417 8435 3451
rect 1501 3349 1535 3383
rect 3525 3349 3559 3383
rect 7113 3349 7147 3383
rect 8677 3349 8711 3383
rect 3065 3145 3099 3179
rect 6830 3145 6864 3179
rect 1777 3077 1811 3111
rect 4353 3077 4387 3111
rect 8953 3077 8987 3111
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 5558 3009 5592 3043
rect 5825 3009 5859 3043
rect 6101 3009 6135 3043
rect 6653 3009 6687 3043
rect 6745 3009 6779 3043
rect 6929 3009 6963 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 7564 3009 7598 3043
rect 6009 2873 6043 2907
rect 1501 2805 1535 2839
rect 4445 2805 4479 2839
rect 7205 2805 7239 2839
rect 8677 2805 8711 2839
rect 9229 2805 9263 2839
rect 4445 2601 4479 2635
rect 5549 2601 5583 2635
rect 6745 2465 6779 2499
rect 7665 2465 7699 2499
rect 1501 2397 1535 2431
rect 1768 2397 1802 2431
rect 3801 2397 3835 2431
rect 5181 2397 5215 2431
rect 5365 2397 5399 2431
rect 6377 2397 6411 2431
rect 7941 2397 7975 2431
rect 9321 2397 9355 2431
rect 3157 2329 3191 2363
rect 3525 2329 3559 2363
rect 4813 2329 4847 2363
rect 6101 2329 6135 2363
rect 6561 2329 6595 2363
rect 7389 2329 7423 2363
rect 2881 2261 2915 2295
rect 5825 2261 5859 2295
rect 8033 2261 8067 2295
rect 9045 2261 9079 2295
<< metal1 >>
rect 1104 10906 10028 10928
rect 1104 10854 2725 10906
rect 2777 10854 2789 10906
rect 2841 10854 2853 10906
rect 2905 10854 2917 10906
rect 2969 10854 2981 10906
rect 3033 10854 4956 10906
rect 5008 10854 5020 10906
rect 5072 10854 5084 10906
rect 5136 10854 5148 10906
rect 5200 10854 5212 10906
rect 5264 10854 7187 10906
rect 7239 10854 7251 10906
rect 7303 10854 7315 10906
rect 7367 10854 7379 10906
rect 7431 10854 7443 10906
rect 7495 10854 9418 10906
rect 9470 10854 9482 10906
rect 9534 10854 9546 10906
rect 9598 10854 9610 10906
rect 9662 10854 9674 10906
rect 9726 10854 10028 10906
rect 1104 10832 10028 10854
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 2240 10724 2268 10755
rect 2590 10752 2596 10804
rect 2648 10792 2654 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2648 10764 2789 10792
rect 2648 10752 2654 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 2777 10755 2835 10761
rect 3050 10752 3056 10804
rect 3108 10752 3114 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 3936 10764 4169 10792
rect 3936 10752 3942 10764
rect 4157 10761 4169 10764
rect 4203 10761 4215 10795
rect 4157 10755 4215 10761
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 5868 10764 6469 10792
rect 5868 10752 5874 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 9306 10752 9312 10804
rect 9364 10752 9370 10804
rect 3068 10724 3096 10752
rect 2240 10696 3096 10724
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2958 10656 2964 10668
rect 2363 10628 2964 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 1780 10588 1808 10619
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 2590 10588 2596 10600
rect 1780 10560 2596 10588
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3068 10464 3096 10619
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 4062 10616 4068 10668
rect 4120 10616 4126 10668
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 4856 10628 6745 10656
rect 4856 10616 4862 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7650 10656 7656 10668
rect 7607 10628 7656 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 8444 10560 8493 10588
rect 8444 10548 8450 10560
rect 8481 10557 8493 10560
rect 8527 10588 8539 10591
rect 9048 10588 9076 10619
rect 8527 10560 9076 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 1486 10412 1492 10464
rect 1544 10412 1550 10464
rect 3050 10412 3056 10464
rect 3108 10412 3114 10464
rect 3234 10412 3240 10464
rect 3292 10412 3298 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7064 10424 7941 10452
rect 7064 10412 7070 10424
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 1104 10362 10028 10384
rect 1104 10310 2065 10362
rect 2117 10310 2129 10362
rect 2181 10310 2193 10362
rect 2245 10310 2257 10362
rect 2309 10310 2321 10362
rect 2373 10310 4296 10362
rect 4348 10310 4360 10362
rect 4412 10310 4424 10362
rect 4476 10310 4488 10362
rect 4540 10310 4552 10362
rect 4604 10310 6527 10362
rect 6579 10310 6591 10362
rect 6643 10310 6655 10362
rect 6707 10310 6719 10362
rect 6771 10310 6783 10362
rect 6835 10310 8758 10362
rect 8810 10310 8822 10362
rect 8874 10310 8886 10362
rect 8938 10310 8950 10362
rect 9002 10310 9014 10362
rect 9066 10310 10028 10362
rect 1104 10288 10028 10310
rect 1302 10208 1308 10260
rect 1360 10248 1366 10260
rect 3329 10251 3387 10257
rect 3329 10248 3341 10251
rect 1360 10220 3341 10248
rect 1360 10208 1366 10220
rect 3329 10217 3341 10220
rect 3375 10217 3387 10251
rect 3329 10211 3387 10217
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3476 10220 3801 10248
rect 3476 10208 3482 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 9585 10251 9643 10257
rect 9585 10217 9597 10251
rect 9631 10248 9643 10251
rect 10318 10248 10324 10260
rect 9631 10220 10324 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 3050 10140 3056 10192
rect 3108 10140 3114 10192
rect 3068 10112 3096 10140
rect 4341 10115 4399 10121
rect 4341 10112 4353 10115
rect 3068 10084 4353 10112
rect 4341 10081 4353 10084
rect 4387 10081 4399 10115
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 4341 10075 4399 10081
rect 6472 10084 7389 10112
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 2498 10044 2504 10056
rect 1719 10016 2504 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5350 10044 5356 10056
rect 4939 10016 5356 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 6472 10044 6500 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 5500 10016 6500 10044
rect 5500 10004 5506 10016
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 1940 9979 1998 9985
rect 1940 9945 1952 9979
rect 1986 9976 1998 9979
rect 2222 9976 2228 9988
rect 1986 9948 2228 9976
rect 1986 9945 1998 9948
rect 1940 9939 1998 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 3237 9979 3295 9985
rect 3237 9976 3249 9979
rect 2424 9948 3249 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2424 9908 2452 9948
rect 3237 9945 3249 9948
rect 3283 9945 3295 9979
rect 4724 9976 4752 10004
rect 4985 9979 5043 9985
rect 4985 9976 4997 9979
rect 4724 9948 4997 9976
rect 3237 9939 3295 9945
rect 4985 9945 4997 9948
rect 5031 9945 5043 9979
rect 4985 9939 5043 9945
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5712 9979 5770 9985
rect 5215 9948 5672 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5644 9920 5672 9948
rect 5712 9945 5724 9979
rect 5758 9976 5770 9979
rect 5810 9976 5816 9988
rect 5758 9948 5816 9976
rect 5758 9945 5770 9948
rect 5712 9939 5770 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 7116 9920 7144 10007
rect 9122 10004 9128 10056
rect 9180 10004 9186 10056
rect 7644 9979 7702 9985
rect 7644 9945 7656 9979
rect 7690 9976 7702 9979
rect 7926 9976 7932 9988
rect 7690 9948 7932 9976
rect 7690 9945 7702 9948
rect 7644 9939 7702 9945
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 9766 9976 9772 9988
rect 9355 9948 9772 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 9766 9936 9772 9948
rect 9824 9936 9830 9988
rect 1627 9880 2452 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 4709 9911 4767 9917
rect 4709 9908 4721 9911
rect 4672 9880 4721 9908
rect 4672 9868 4678 9880
rect 4709 9877 4721 9880
rect 4755 9877 4767 9911
rect 4709 9871 4767 9877
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 5534 9908 5540 9920
rect 5399 9880 5540 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 6825 9911 6883 9917
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 7006 9908 7012 9920
rect 6871 9880 7012 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7098 9868 7104 9920
rect 7156 9868 7162 9920
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 8018 9908 8024 9920
rect 7331 9880 8024 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8444 9880 8769 9908
rect 8444 9868 8450 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 8938 9868 8944 9920
rect 8996 9868 9002 9920
rect 1104 9818 10028 9840
rect 1104 9766 2725 9818
rect 2777 9766 2789 9818
rect 2841 9766 2853 9818
rect 2905 9766 2917 9818
rect 2969 9766 2981 9818
rect 3033 9766 4956 9818
rect 5008 9766 5020 9818
rect 5072 9766 5084 9818
rect 5136 9766 5148 9818
rect 5200 9766 5212 9818
rect 5264 9766 7187 9818
rect 7239 9766 7251 9818
rect 7303 9766 7315 9818
rect 7367 9766 7379 9818
rect 7431 9766 7443 9818
rect 7495 9766 9418 9818
rect 9470 9766 9482 9818
rect 9534 9766 9546 9818
rect 9598 9766 9610 9818
rect 9662 9766 9674 9818
rect 9726 9766 10028 9818
rect 1104 9744 10028 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 1452 9676 2176 9704
rect 1452 9664 1458 9676
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 2148 9636 2176 9676
rect 2222 9664 2228 9716
rect 2280 9664 2286 9716
rect 3605 9707 3663 9713
rect 2332 9676 3556 9704
rect 2332 9636 2360 9676
rect 2148 9608 2360 9636
rect 3528 9636 3556 9676
rect 3605 9673 3617 9707
rect 3651 9704 3663 9707
rect 4062 9704 4068 9716
rect 3651 9676 4068 9704
rect 3651 9673 3663 9676
rect 3605 9667 3663 9673
rect 4062 9664 4068 9676
rect 4120 9664 4126 9716
rect 5534 9664 5540 9716
rect 5592 9664 5598 9716
rect 5626 9664 5632 9716
rect 5684 9664 5690 9716
rect 5810 9664 5816 9716
rect 5868 9664 5874 9716
rect 3528 9608 4200 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 3234 9568 3240 9580
rect 2455 9540 3240 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 1964 9432 1992 9531
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3467 9540 4108 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3234 9432 3240 9444
rect 1964 9404 3240 9432
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 4080 9376 4108 9540
rect 4172 9376 4200 9608
rect 4614 9528 4620 9580
rect 4672 9568 4678 9580
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 4672 9540 4721 9568
rect 4672 9528 4678 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 4709 9531 4767 9537
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4856 9540 5089 9568
rect 4856 9528 4862 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9537 5503 9571
rect 5552 9568 5580 9664
rect 5644 9636 5672 9664
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 5644 9608 6377 9636
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 7285 9639 7343 9645
rect 7285 9605 7297 9639
rect 7331 9636 7343 9639
rect 8386 9636 8392 9648
rect 7331 9608 8392 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 8564 9639 8622 9645
rect 8564 9605 8576 9639
rect 8610 9636 8622 9639
rect 8938 9636 8944 9648
rect 8610 9608 8944 9636
rect 8610 9605 8622 9608
rect 8564 9599 8622 9605
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5552 9540 5641 9568
rect 5445 9531 5503 9537
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 7098 9568 7104 9580
rect 5629 9531 5687 9537
rect 6932 9540 7104 9568
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5460 9432 5488 9531
rect 6932 9432 6960 9540
rect 7098 9528 7104 9540
rect 7156 9568 7162 9580
rect 7469 9571 7527 9577
rect 7469 9568 7481 9571
rect 7156 9540 7481 9568
rect 7156 9528 7162 9540
rect 7469 9537 7481 9540
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7650 9500 7656 9512
rect 7064 9472 7656 9500
rect 7064 9460 7070 9472
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8294 9460 8300 9512
rect 8352 9460 8358 9512
rect 5123 9404 6960 9432
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 6932 9376 6960 9404
rect 9677 9435 9735 9441
rect 9677 9401 9689 9435
rect 9723 9432 9735 9435
rect 9766 9432 9772 9444
rect 9723 9404 9772 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 1820 9336 2513 9364
rect 1820 9324 1826 9336
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 2501 9327 2559 9333
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 4062 9364 4068 9376
rect 2740 9336 4068 9364
rect 2740 9324 2746 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4706 9364 4712 9376
rect 4212 9336 4712 9364
rect 4212 9324 4218 9336
rect 4706 9324 4712 9336
rect 4764 9364 4770 9376
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 4764 9336 5365 9364
rect 4764 9324 4770 9336
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5353 9327 5411 9333
rect 6914 9324 6920 9376
rect 6972 9324 6978 9376
rect 7098 9324 7104 9376
rect 7156 9324 7162 9376
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8202 9364 8208 9376
rect 8067 9336 8208 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8202 9324 8208 9336
rect 8260 9324 8266 9376
rect 1104 9274 10028 9296
rect 1104 9222 2065 9274
rect 2117 9222 2129 9274
rect 2181 9222 2193 9274
rect 2245 9222 2257 9274
rect 2309 9222 2321 9274
rect 2373 9222 4296 9274
rect 4348 9222 4360 9274
rect 4412 9222 4424 9274
rect 4476 9222 4488 9274
rect 4540 9222 4552 9274
rect 4604 9222 6527 9274
rect 6579 9222 6591 9274
rect 6643 9222 6655 9274
rect 6707 9222 6719 9274
rect 6771 9222 6783 9274
rect 6835 9222 8758 9274
rect 8810 9222 8822 9274
rect 8874 9222 8886 9274
rect 8938 9222 8950 9274
rect 9002 9222 9014 9274
rect 9066 9222 10028 9274
rect 1104 9200 10028 9222
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 3108 9132 3341 9160
rect 3108 9120 3114 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 7561 9163 7619 9169
rect 4120 9132 7144 9160
rect 4120 9120 4126 9132
rect 3234 9052 3240 9104
rect 3292 9092 3298 9104
rect 5350 9092 5356 9104
rect 3292 9064 5356 9092
rect 3292 9052 3298 9064
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 7116 9092 7144 9132
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 7834 9160 7840 9172
rect 7607 9132 7840 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 7926 9120 7932 9172
rect 7984 9120 7990 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8205 9163 8263 9169
rect 8205 9160 8217 9163
rect 8168 9132 8217 9160
rect 8168 9120 8174 9132
rect 8205 9129 8217 9132
rect 8251 9129 8263 9163
rect 8205 9123 8263 9129
rect 7116 9064 8432 9092
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 9024 1639 9027
rect 2498 9024 2504 9036
rect 1627 8996 2504 9024
rect 1627 8993 1639 8996
rect 1581 8987 1639 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 4614 9024 4620 9036
rect 3844 8996 4620 9024
rect 3844 8984 3850 8996
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 8294 9024 8300 9036
rect 5828 8996 8300 9024
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 3651 8928 4108 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 1854 8848 1860 8900
rect 1912 8848 1918 8900
rect 3513 8891 3571 8897
rect 3513 8888 3525 8891
rect 3082 8860 3525 8888
rect 3513 8857 3525 8860
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 4080 8832 4108 8928
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5442 8956 5448 8968
rect 4856 8928 5448 8956
rect 4856 8916 4862 8928
rect 5442 8916 5448 8928
rect 5500 8956 5506 8968
rect 5828 8965 5856 8996
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8404 9024 8432 9064
rect 8570 9024 8576 9036
rect 8404 8996 8576 9024
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5500 8928 5825 8956
rect 5500 8916 5506 8928
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 6086 8848 6092 8900
rect 6144 8848 6150 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7314 8860 7757 8888
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2682 8820 2688 8832
rect 2280 8792 2688 8820
rect 2280 8780 2286 8792
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 7852 8820 7880 8919
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8404 8965 8432 8996
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 8113 8959 8171 8965
rect 8113 8956 8125 8959
rect 8076 8928 8125 8956
rect 8076 8916 8082 8928
rect 8113 8925 8125 8928
rect 8159 8925 8171 8959
rect 8113 8919 8171 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 7926 8848 7932 8900
rect 7984 8888 7990 8900
rect 8496 8888 8524 8919
rect 9674 8888 9680 8900
rect 7984 8860 8524 8888
rect 8680 8860 9680 8888
rect 7984 8848 7990 8860
rect 8478 8820 8484 8832
rect 4120 8792 8484 8820
rect 4120 8780 4126 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8680 8829 8708 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 8665 8823 8723 8829
rect 8665 8789 8677 8823
rect 8711 8789 8723 8823
rect 8665 8783 8723 8789
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 1104 8730 10028 8752
rect 1104 8678 2725 8730
rect 2777 8678 2789 8730
rect 2841 8678 2853 8730
rect 2905 8678 2917 8730
rect 2969 8678 2981 8730
rect 3033 8678 4956 8730
rect 5008 8678 5020 8730
rect 5072 8678 5084 8730
rect 5136 8678 5148 8730
rect 5200 8678 5212 8730
rect 5264 8678 7187 8730
rect 7239 8678 7251 8730
rect 7303 8678 7315 8730
rect 7367 8678 7379 8730
rect 7431 8678 7443 8730
rect 7495 8678 9418 8730
rect 9470 8678 9482 8730
rect 9534 8678 9546 8730
rect 9598 8678 9610 8730
rect 9662 8678 9674 8730
rect 9726 8678 10028 8730
rect 1104 8656 10028 8678
rect 1762 8576 1768 8628
rect 1820 8576 1826 8628
rect 1854 8576 1860 8628
rect 1912 8576 1918 8628
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2317 8619 2375 8625
rect 2317 8616 2329 8619
rect 2280 8588 2329 8616
rect 2280 8576 2286 8588
rect 2317 8585 2329 8588
rect 2363 8585 2375 8619
rect 2317 8579 2375 8585
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 1780 8480 1808 8576
rect 1627 8452 1808 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 1872 8412 1900 8576
rect 2332 8548 2360 8579
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 3050 8616 3056 8628
rect 2556 8588 3056 8616
rect 2556 8576 2562 8588
rect 2332 8520 2544 8548
rect 2516 8492 2544 8520
rect 2406 8440 2412 8492
rect 2464 8440 2470 8492
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2700 8489 2728 8588
rect 3050 8576 3056 8588
rect 3108 8616 3114 8628
rect 4798 8616 4804 8628
rect 3108 8588 4804 8616
rect 3108 8576 3114 8588
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 7834 8616 7840 8628
rect 5408 8588 7840 8616
rect 5408 8576 5414 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 3970 8508 3976 8560
rect 4028 8508 4034 8560
rect 4706 8508 4712 8560
rect 4764 8508 4770 8560
rect 4816 8489 4844 8576
rect 5074 8489 5080 8492
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 5068 8443 5080 8489
rect 1949 8415 2007 8421
rect 1949 8412 1961 8415
rect 1872 8384 1961 8412
rect 1949 8381 1961 8384
rect 1995 8381 2007 8415
rect 2608 8412 2636 8443
rect 5074 8440 5080 8443
rect 5132 8440 5138 8492
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9048 8480 9076 8576
rect 8895 8452 9076 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9364 8452 9505 8480
rect 9364 8440 9370 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 2608 8384 2973 8412
rect 1949 8375 2007 8381
rect 2961 8381 2973 8384
rect 3007 8412 3019 8415
rect 3326 8412 3332 8424
rect 3007 8384 3332 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 9122 8372 9128 8424
rect 9180 8372 9186 8424
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 9140 8344 9168 8372
rect 9079 8316 9168 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 6196 8276 6224 8307
rect 7926 8276 7932 8288
rect 6196 8248 7932 8276
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 1104 8186 10028 8208
rect 1104 8134 2065 8186
rect 2117 8134 2129 8186
rect 2181 8134 2193 8186
rect 2245 8134 2257 8186
rect 2309 8134 2321 8186
rect 2373 8134 4296 8186
rect 4348 8134 4360 8186
rect 4412 8134 4424 8186
rect 4476 8134 4488 8186
rect 4540 8134 4552 8186
rect 4604 8134 6527 8186
rect 6579 8134 6591 8186
rect 6643 8134 6655 8186
rect 6707 8134 6719 8186
rect 6771 8134 6783 8186
rect 6835 8134 8758 8186
rect 8810 8134 8822 8186
rect 8874 8134 8886 8186
rect 8938 8134 8950 8186
rect 9002 8134 9014 8186
rect 9066 8134 10028 8186
rect 1104 8112 10028 8134
rect 934 8032 940 8084
rect 992 8072 998 8084
rect 1489 8075 1547 8081
rect 1489 8072 1501 8075
rect 992 8044 1501 8072
rect 992 8032 998 8044
rect 1489 8041 1501 8044
rect 1535 8041 1547 8075
rect 1489 8035 1547 8041
rect 3326 8032 3332 8084
rect 3384 8032 3390 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 3970 8072 3976 8084
rect 3927 8044 3976 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4985 8075 5043 8081
rect 4985 8041 4997 8075
rect 5031 8072 5043 8075
rect 5074 8072 5080 8084
rect 5031 8044 5080 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6144 8044 6193 8072
rect 6144 8032 6150 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 7742 8004 7748 8016
rect 6104 7976 7748 8004
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 2406 7936 2412 7948
rect 2087 7908 2412 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 2056 7868 2084 7899
rect 2406 7896 2412 7908
rect 2464 7936 2470 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 2464 7908 3004 7936
rect 2464 7896 2470 7908
rect 1811 7840 2084 7868
rect 2133 7871 2191 7877
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 2179 7840 2452 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2424 7744 2452 7840
rect 2590 7828 2596 7880
rect 2648 7868 2654 7880
rect 2976 7877 3004 7908
rect 3436 7908 4077 7936
rect 3436 7877 3464 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4065 7899 4123 7905
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 2961 7871 3019 7877
rect 2648 7840 2820 7868
rect 2648 7828 2654 7840
rect 2792 7809 2820 7840
rect 2961 7837 2973 7871
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3568 7840 3985 7868
rect 3568 7828 3574 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3988 7800 4016 7831
rect 4798 7828 4804 7880
rect 4856 7828 4862 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6104 7877 6132 7976
rect 6932 7945 6960 7976
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 6917 7939 6975 7945
rect 6288 7908 6868 7936
rect 6288 7877 6316 7908
rect 6840 7880 6868 7908
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 6917 7899 6975 7905
rect 7006 7896 7012 7948
rect 7064 7896 7070 7948
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5960 7840 6101 7868
rect 5960 7828 5966 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6420 7840 6745 7868
rect 6420 7828 6426 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7837 7159 7871
rect 7208 7868 7236 7896
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 7208 7840 7297 7868
rect 7101 7831 7159 7837
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 4062 7800 4068 7812
rect 2823 7772 3464 7800
rect 3988 7772 4068 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 3436 7744 3464 7772
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 7116 7800 7144 7831
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 6104 7772 7144 7800
rect 7208 7772 9321 7800
rect 6104 7744 6132 7772
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 3142 7692 3148 7744
rect 3200 7692 3206 7744
rect 3418 7692 3424 7744
rect 3476 7692 3482 7744
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6328 7704 6561 7732
rect 6328 7692 6334 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6549 7695 6607 7701
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7208 7732 7236 7772
rect 9309 7769 9321 7772
rect 9355 7800 9367 7803
rect 9355 7772 10088 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 7064 7704 7236 7732
rect 8297 7735 8355 7741
rect 7064 7692 7070 7704
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8386 7732 8392 7744
rect 8343 7704 8392 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9585 7735 9643 7741
rect 9585 7701 9597 7735
rect 9631 7732 9643 7735
rect 9950 7732 9956 7744
rect 9631 7704 9956 7732
rect 9631 7701 9643 7704
rect 9585 7695 9643 7701
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 1104 7642 10028 7664
rect 1104 7590 2725 7642
rect 2777 7590 2789 7642
rect 2841 7590 2853 7642
rect 2905 7590 2917 7642
rect 2969 7590 2981 7642
rect 3033 7590 4956 7642
rect 5008 7590 5020 7642
rect 5072 7590 5084 7642
rect 5136 7590 5148 7642
rect 5200 7590 5212 7642
rect 5264 7590 7187 7642
rect 7239 7590 7251 7642
rect 7303 7590 7315 7642
rect 7367 7590 7379 7642
rect 7431 7590 7443 7642
rect 7495 7590 9418 7642
rect 9470 7590 9482 7642
rect 9534 7590 9546 7642
rect 9598 7590 9610 7642
rect 9662 7590 9674 7642
rect 9726 7590 10028 7642
rect 1104 7568 10028 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3050 7528 3056 7540
rect 2915 7500 3056 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3142 7488 3148 7540
rect 3200 7488 3206 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 5077 7531 5135 7537
rect 5077 7528 5089 7531
rect 4856 7500 5089 7528
rect 4856 7488 4862 7500
rect 5077 7497 5089 7500
rect 5123 7497 5135 7531
rect 5077 7491 5135 7497
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 7006 7528 7012 7540
rect 6687 7500 7012 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 9677 7531 9735 7537
rect 9677 7497 9689 7531
rect 9723 7528 9735 7531
rect 10060 7528 10088 7772
rect 9723 7500 10088 7528
rect 9723 7497 9735 7500
rect 9677 7491 9735 7497
rect 3160 7324 3188 7488
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 4614 7460 4620 7472
rect 4387 7432 4620 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 4614 7420 4620 7432
rect 4672 7420 4678 7472
rect 5261 7463 5319 7469
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 5350 7460 5356 7472
rect 5307 7432 5356 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 5350 7420 5356 7432
rect 5408 7460 5414 7472
rect 7466 7460 7472 7472
rect 5408 7432 7472 7460
rect 5408 7420 5414 7432
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4212 7364 4905 7392
rect 4212 7352 4218 7364
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 4617 7327 4675 7333
rect 4617 7324 4629 7327
rect 3160 7296 4629 7324
rect 4617 7293 4629 7296
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4706 7284 4712 7336
rect 4764 7284 4770 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4908 7324 4936 7355
rect 5442 7352 5448 7404
rect 5500 7352 5506 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 7392 7401 7420 7432
rect 7466 7420 7472 7432
rect 7524 7460 7530 7472
rect 7944 7460 7972 7488
rect 7524 7432 7972 7460
rect 8404 7460 8432 7488
rect 8542 7463 8600 7469
rect 8542 7460 8554 7463
rect 8404 7432 8554 7460
rect 7524 7420 7530 7432
rect 8542 7429 8554 7432
rect 8588 7429 8600 7463
rect 8542 7423 8600 7429
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6420 7364 6745 7392
rect 6420 7352 6426 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7650 7352 7656 7404
rect 7708 7352 7714 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8018 7392 8024 7404
rect 7975 7364 8024 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 4908 7296 6469 7324
rect 4801 7287 4859 7293
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 4816 7256 4844 7287
rect 7558 7284 7564 7336
rect 7616 7284 7622 7336
rect 7760 7324 7788 7355
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 7668 7296 7788 7324
rect 8220 7324 8248 7355
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8404 7324 8432 7352
rect 8220 7296 8432 7324
rect 7668 7268 7696 7296
rect 4816 7228 5028 7256
rect 5000 7200 5028 7228
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 7650 7256 7656 7268
rect 6880 7228 7656 7256
rect 6880 7216 6886 7228
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4798 7188 4804 7200
rect 4479 7160 4804 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 4982 7148 4988 7200
rect 5040 7148 5046 7200
rect 7098 7148 7104 7200
rect 7156 7148 7162 7200
rect 7190 7148 7196 7200
rect 7248 7148 7254 7200
rect 8113 7191 8171 7197
rect 8113 7157 8125 7191
rect 8159 7188 8171 7191
rect 8202 7188 8208 7200
rect 8159 7160 8208 7188
rect 8159 7157 8171 7160
rect 8113 7151 8171 7157
rect 8202 7148 8208 7160
rect 8260 7148 8266 7200
rect 1104 7098 10028 7120
rect 1104 7046 2065 7098
rect 2117 7046 2129 7098
rect 2181 7046 2193 7098
rect 2245 7046 2257 7098
rect 2309 7046 2321 7098
rect 2373 7046 4296 7098
rect 4348 7046 4360 7098
rect 4412 7046 4424 7098
rect 4476 7046 4488 7098
rect 4540 7046 4552 7098
rect 4604 7046 6527 7098
rect 6579 7046 6591 7098
rect 6643 7046 6655 7098
rect 6707 7046 6719 7098
rect 6771 7046 6783 7098
rect 6835 7046 8758 7098
rect 8810 7046 8822 7098
rect 8874 7046 8886 7098
rect 8938 7046 8950 7098
rect 9002 7046 9014 7098
rect 9066 7046 10028 7098
rect 1104 7024 10028 7046
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 3786 6984 3792 6996
rect 2464 6956 3792 6984
rect 2464 6944 2470 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4246 6944 4252 6996
rect 4304 6984 4310 6996
rect 4890 6984 4896 6996
rect 4304 6956 4896 6984
rect 4304 6944 4310 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 7098 6944 7104 6996
rect 7156 6944 7162 6996
rect 7742 6944 7748 6996
rect 7800 6944 7806 6996
rect 8018 6944 8024 6996
rect 8076 6944 8082 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8444 6956 8953 6984
rect 8444 6944 8450 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 4672 6888 5580 6916
rect 4672 6876 4678 6888
rect 2777 6851 2835 6857
rect 2777 6848 2789 6851
rect 2240 6820 2789 6848
rect 1670 6740 1676 6792
rect 1728 6780 1734 6792
rect 1946 6780 1952 6792
rect 1728 6752 1952 6780
rect 1728 6740 1734 6752
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6782 2191 6783
rect 2240 6782 2268 6820
rect 2777 6817 2789 6820
rect 2823 6817 2835 6851
rect 3326 6848 3332 6860
rect 2777 6811 2835 6817
rect 3160 6820 3332 6848
rect 2179 6754 2268 6782
rect 2179 6749 2191 6754
rect 2133 6743 2191 6749
rect 2682 6740 2688 6792
rect 2740 6740 2746 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1397 6715 1455 6721
rect 1397 6712 1409 6715
rect 992 6684 1409 6712
rect 992 6672 998 6684
rect 1397 6681 1409 6684
rect 1443 6681 1455 6715
rect 1397 6675 1455 6681
rect 1765 6715 1823 6721
rect 1765 6681 1777 6715
rect 1811 6681 1823 6715
rect 2593 6715 2651 6721
rect 1765 6675 1823 6681
rect 2148 6684 2360 6712
rect 1780 6644 1808 6675
rect 2148 6644 2176 6684
rect 1780 6616 2176 6644
rect 2222 6604 2228 6656
rect 2280 6604 2286 6656
rect 2332 6644 2360 6684
rect 2593 6681 2605 6715
rect 2639 6681 2651 6715
rect 2884 6712 2912 6743
rect 3050 6740 3056 6792
rect 3108 6740 3114 6792
rect 3160 6789 3188 6820
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 4154 6848 4160 6860
rect 3559 6820 4160 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 5552 6848 5580 6888
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 5552 6820 6469 6848
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6733 6851 6791 6857
rect 6733 6817 6745 6851
rect 6779 6848 6791 6851
rect 6914 6848 6920 6860
rect 6779 6820 6920 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7116 6848 7144 6944
rect 8680 6888 9168 6916
rect 7055 6820 7144 6848
rect 7484 6820 7972 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7484 6792 7512 6820
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3651 6752 4108 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 2884 6684 3801 6712
rect 2593 6675 2651 6681
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 2393 6647 2451 6653
rect 2393 6644 2405 6647
rect 2332 6616 2405 6644
rect 2393 6613 2405 6616
rect 2439 6644 2451 6647
rect 2498 6644 2504 6656
rect 2439 6616 2504 6644
rect 2439 6613 2451 6616
rect 2393 6607 2451 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2608 6644 2636 6675
rect 3878 6644 3884 6656
rect 2608 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4080 6644 4108 6752
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4488 6752 4629 6780
rect 4488 6740 4494 6752
rect 4617 6749 4629 6752
rect 4663 6780 4675 6783
rect 4982 6780 4988 6792
rect 4663 6752 4988 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 6270 6740 6276 6792
rect 6328 6780 6334 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6328 6752 7113 6780
rect 6328 6740 6334 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7944 6780 7972 6820
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 8680 6848 8708 6888
rect 8076 6820 8708 6848
rect 8076 6808 8082 6820
rect 8754 6808 8760 6860
rect 8812 6808 8818 6860
rect 9140 6857 9168 6888
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9217 6783 9275 6789
rect 9048 6780 9168 6782
rect 9217 6780 9229 6783
rect 7944 6754 9229 6780
rect 7944 6752 9076 6754
rect 9140 6752 9229 6754
rect 7837 6743 7895 6749
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 4893 6715 4951 6721
rect 4893 6712 4905 6715
rect 4212 6684 4905 6712
rect 4212 6672 4218 6684
rect 4893 6681 4905 6684
rect 4939 6681 4951 6715
rect 5000 6712 5028 6740
rect 7558 6712 7564 6724
rect 5000 6684 7564 6712
rect 4893 6675 4951 6681
rect 7558 6672 7564 6684
rect 7616 6672 7622 6724
rect 7852 6712 7880 6743
rect 8113 6715 8171 6721
rect 8113 6712 8125 6715
rect 7852 6684 8125 6712
rect 8113 6681 8125 6684
rect 8159 6681 8171 6715
rect 8113 6675 8171 6681
rect 9585 6715 9643 6721
rect 9585 6681 9597 6715
rect 9631 6681 9643 6715
rect 9585 6675 9643 6681
rect 4522 6644 4528 6656
rect 4080 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 5442 6644 5448 6656
rect 4755 6616 5448 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 8128 6644 8156 6675
rect 9600 6644 9628 6675
rect 8128 6616 9628 6644
rect 1104 6554 10028 6576
rect 1104 6502 2725 6554
rect 2777 6502 2789 6554
rect 2841 6502 2853 6554
rect 2905 6502 2917 6554
rect 2969 6502 2981 6554
rect 3033 6502 4956 6554
rect 5008 6502 5020 6554
rect 5072 6502 5084 6554
rect 5136 6502 5148 6554
rect 5200 6502 5212 6554
rect 5264 6502 7187 6554
rect 7239 6502 7251 6554
rect 7303 6502 7315 6554
rect 7367 6502 7379 6554
rect 7431 6502 7443 6554
rect 7495 6502 9418 6554
rect 9470 6502 9482 6554
rect 9534 6502 9546 6554
rect 9598 6502 9610 6554
rect 9662 6502 9674 6554
rect 9726 6502 10028 6554
rect 1104 6480 10028 6502
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2556 6412 3157 6440
rect 2556 6400 2562 6412
rect 3145 6409 3157 6412
rect 3191 6440 3203 6443
rect 4338 6440 4344 6452
rect 3191 6412 4344 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 4706 6440 4712 6452
rect 4580 6412 4712 6440
rect 4580 6400 4586 6412
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 6917 6443 6975 6449
rect 6917 6440 6929 6443
rect 6420 6412 6929 6440
rect 6420 6400 6426 6412
rect 6917 6409 6929 6412
rect 6963 6409 6975 6443
rect 6917 6403 6975 6409
rect 7006 6400 7012 6452
rect 7064 6400 7070 6452
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 8110 6440 8116 6452
rect 7883 6412 8116 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9306 6440 9312 6452
rect 8812 6412 9312 6440
rect 8812 6400 8818 6412
rect 9306 6400 9312 6412
rect 9364 6440 9370 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9364 6412 9505 6440
rect 9364 6400 9370 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 1673 6375 1731 6381
rect 1673 6341 1685 6375
rect 1719 6372 1731 6375
rect 2056 6372 2084 6400
rect 3050 6372 3056 6384
rect 1719 6344 2084 6372
rect 2898 6344 3056 6372
rect 1719 6341 1731 6344
rect 1673 6335 1731 6341
rect 3050 6332 3056 6344
rect 3108 6332 3114 6384
rect 3602 6332 3608 6384
rect 3660 6332 3666 6384
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 4724 6372 4752 6400
rect 3844 6344 4200 6372
rect 4724 6344 5212 6372
rect 3844 6332 3850 6344
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3467 6276 3832 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 3237 6239 3295 6245
rect 1443 6208 2774 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2746 6168 2774 6208
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3510 6236 3516 6248
rect 3283 6208 3516 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 3804 6236 3832 6276
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 4172 6313 4200 6344
rect 3973 6307 4031 6313
rect 3973 6304 3985 6307
rect 3936 6276 3985 6304
rect 3936 6264 3942 6276
rect 3973 6273 3985 6276
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4157 6307 4215 6313
rect 4338 6308 4344 6316
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4280 6304 4344 6308
rect 4203 6280 4344 6304
rect 4203 6276 4308 6280
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 3988 6236 4016 6267
rect 4338 6264 4344 6280
rect 4396 6264 4402 6316
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6302 4491 6307
rect 4522 6302 4528 6316
rect 4479 6274 4528 6302
rect 4479 6273 4491 6274
rect 4433 6267 4491 6273
rect 4522 6264 4528 6274
rect 4580 6264 4586 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 5074 6304 5080 6316
rect 4764 6276 5080 6304
rect 4764 6264 4770 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5184 6313 5212 6344
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 7024 6304 7052 6400
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 7024 6276 7113 6304
rect 6917 6267 6975 6273
rect 7101 6273 7113 6276
rect 7147 6304 7159 6307
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7147 6276 7481 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7576 6304 7604 6400
rect 8202 6332 8208 6384
rect 8260 6332 8266 6384
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7576 6276 7665 6304
rect 7469 6267 7527 6273
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 8220 6304 8248 6332
rect 8369 6307 8427 6313
rect 8369 6304 8381 6307
rect 8220 6276 8381 6304
rect 7653 6267 7711 6273
rect 8369 6273 8381 6276
rect 8415 6273 8427 6307
rect 8369 6267 8427 6273
rect 4246 6236 4252 6248
rect 3804 6208 3924 6236
rect 3988 6208 4252 6236
rect 3620 6168 3648 6196
rect 2746 6140 3648 6168
rect 3896 6168 3924 6208
rect 4246 6196 4252 6208
rect 4304 6236 4310 6248
rect 4801 6239 4859 6245
rect 4304 6208 4752 6236
rect 4304 6196 4310 6208
rect 4430 6168 4436 6180
rect 3896 6140 4436 6168
rect 3896 6109 3924 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 4724 6168 4752 6208
rect 4801 6205 4813 6239
rect 4847 6236 4859 6239
rect 4890 6236 4896 6248
rect 4847 6208 4896 6236
rect 4847 6205 4859 6208
rect 4801 6199 4859 6205
rect 4890 6196 4896 6208
rect 4948 6236 4954 6248
rect 5368 6236 5396 6264
rect 4948 6208 5396 6236
rect 4948 6196 4954 6208
rect 5442 6196 5448 6248
rect 5500 6196 5506 6248
rect 6932 6236 6960 6267
rect 7834 6236 7840 6248
rect 6932 6208 7840 6236
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 7926 6196 7932 6248
rect 7984 6236 7990 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7984 6208 8125 6236
rect 7984 6196 7990 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 7006 6168 7012 6180
rect 4724 6140 7012 6168
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6069 3939 6103
rect 3881 6063 3939 6069
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 4028 6072 4261 6100
rect 4028 6060 4034 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4706 6100 4712 6112
rect 4396 6072 4712 6100
rect 4396 6060 4402 6072
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 4982 6060 4988 6112
rect 5040 6060 5046 6112
rect 5258 6060 5264 6112
rect 5316 6060 5322 6112
rect 5718 6060 5724 6112
rect 5776 6060 5782 6112
rect 1104 6010 10028 6032
rect 1104 5958 2065 6010
rect 2117 5958 2129 6010
rect 2181 5958 2193 6010
rect 2245 5958 2257 6010
rect 2309 5958 2321 6010
rect 2373 5958 4296 6010
rect 4348 5958 4360 6010
rect 4412 5958 4424 6010
rect 4476 5958 4488 6010
rect 4540 5958 4552 6010
rect 4604 5958 6527 6010
rect 6579 5958 6591 6010
rect 6643 5958 6655 6010
rect 6707 5958 6719 6010
rect 6771 5958 6783 6010
rect 6835 5958 8758 6010
rect 8810 5958 8822 6010
rect 8874 5958 8886 6010
rect 8938 5958 8950 6010
rect 9002 5958 9014 6010
rect 9066 5958 10028 6010
rect 1104 5936 10028 5958
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 3418 5896 3424 5908
rect 2271 5868 3424 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 4249 5899 4307 5905
rect 4249 5865 4261 5899
rect 4295 5865 4307 5899
rect 4249 5859 4307 5865
rect 3988 5760 4016 5856
rect 3528 5732 4016 5760
rect 4264 5760 4292 5859
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 4985 5899 5043 5905
rect 4985 5896 4997 5899
rect 4948 5868 4997 5896
rect 4948 5856 4954 5868
rect 4985 5865 4997 5868
rect 5031 5865 5043 5899
rect 4985 5859 5043 5865
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 5258 5896 5264 5908
rect 5215 5868 5264 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 6641 5899 6699 5905
rect 6641 5865 6653 5899
rect 6687 5865 6699 5899
rect 6641 5859 6699 5865
rect 6656 5828 6684 5859
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8018 5896 8024 5908
rect 7892 5868 8024 5896
rect 7892 5856 7898 5868
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 9306 5828 9312 5840
rect 6656 5800 9312 5828
rect 9306 5788 9312 5800
rect 9364 5828 9370 5840
rect 9364 5800 9536 5828
rect 9364 5788 9370 5800
rect 9508 5769 9536 5800
rect 7285 5763 7343 5769
rect 4264 5732 7144 5760
rect 3349 5695 3407 5701
rect 3349 5661 3361 5695
rect 3395 5692 3407 5695
rect 3528 5692 3556 5732
rect 3395 5664 3556 5692
rect 3395 5661 3407 5664
rect 3349 5655 3407 5661
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 3878 5692 3884 5704
rect 3660 5664 3884 5692
rect 3660 5652 3666 5664
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4172 5664 4936 5692
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 1765 5627 1823 5633
rect 1765 5624 1777 5627
rect 1452 5596 1777 5624
rect 1452 5584 1458 5596
rect 1765 5593 1777 5596
rect 1811 5593 1823 5627
rect 1765 5587 1823 5593
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 4065 5627 4123 5633
rect 4065 5624 4077 5627
rect 3568 5596 4077 5624
rect 3568 5584 3574 5596
rect 4065 5593 4077 5596
rect 4111 5593 4123 5627
rect 4065 5587 4123 5593
rect 4172 5568 4200 5664
rect 4801 5627 4859 5633
rect 4801 5593 4813 5627
rect 4847 5593 4859 5627
rect 4908 5624 4936 5664
rect 5902 5652 5908 5704
rect 5960 5652 5966 5704
rect 6012 5701 6040 5732
rect 5997 5695 6055 5701
rect 5997 5661 6009 5695
rect 6043 5661 6055 5695
rect 5997 5655 6055 5661
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6411 5664 6500 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 4982 5624 4988 5636
rect 5040 5633 5046 5636
rect 5040 5627 5059 5633
rect 4908 5596 4988 5624
rect 4801 5587 4859 5593
rect 1854 5516 1860 5568
rect 1912 5516 1918 5568
rect 4154 5516 4160 5568
rect 4212 5516 4218 5568
rect 4246 5516 4252 5568
rect 4304 5565 4310 5568
rect 4304 5559 4323 5565
rect 4311 5525 4323 5559
rect 4304 5519 4323 5525
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4706 5556 4712 5568
rect 4479 5528 4712 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4304 5516 4310 5519
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 4816 5556 4844 5587
rect 4982 5584 4988 5596
rect 5047 5624 5059 5627
rect 6089 5627 6147 5633
rect 6089 5624 6101 5627
rect 5047 5596 6101 5624
rect 5047 5593 5059 5596
rect 5040 5587 5059 5593
rect 6089 5593 6101 5596
rect 6135 5593 6147 5627
rect 6089 5587 6147 5593
rect 5040 5584 5046 5587
rect 5166 5556 5172 5568
rect 4816 5528 5172 5556
rect 5166 5516 5172 5528
rect 5224 5556 5230 5568
rect 5350 5556 5356 5568
rect 5224 5528 5356 5556
rect 5224 5516 5230 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6472 5565 6500 5664
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6604 5664 7021 5692
rect 6604 5652 6610 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7116 5692 7144 5732
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 7331 5732 8953 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7116 5664 7481 5692
rect 7009 5655 7067 5661
rect 7469 5661 7481 5664
rect 7515 5692 7527 5695
rect 7558 5692 7564 5704
rect 7515 5664 7564 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7699 5664 7849 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 5721 5559 5779 5565
rect 5721 5556 5733 5559
rect 5684 5528 5733 5556
rect 5684 5516 5690 5528
rect 5721 5525 5733 5528
rect 5767 5525 5779 5559
rect 5721 5519 5779 5525
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5525 6515 5559
rect 6457 5519 6515 5525
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6822 5556 6828 5568
rect 6687 5528 6828 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6822 5516 6828 5528
rect 6880 5556 6886 5568
rect 7006 5556 7012 5568
rect 6880 5528 7012 5556
rect 6880 5516 6886 5528
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 8018 5516 8024 5568
rect 8076 5516 8082 5568
rect 1104 5466 10028 5488
rect 1104 5414 2725 5466
rect 2777 5414 2789 5466
rect 2841 5414 2853 5466
rect 2905 5414 2917 5466
rect 2969 5414 2981 5466
rect 3033 5414 4956 5466
rect 5008 5414 5020 5466
rect 5072 5414 5084 5466
rect 5136 5414 5148 5466
rect 5200 5414 5212 5466
rect 5264 5414 7187 5466
rect 7239 5414 7251 5466
rect 7303 5414 7315 5466
rect 7367 5414 7379 5466
rect 7431 5414 7443 5466
rect 7495 5414 9418 5466
rect 9470 5414 9482 5466
rect 9534 5414 9546 5466
rect 9598 5414 9610 5466
rect 9662 5414 9674 5466
rect 9726 5414 10028 5466
rect 1104 5392 10028 5414
rect 4246 5312 4252 5364
rect 4304 5352 4310 5364
rect 4341 5355 4399 5361
rect 4341 5352 4353 5355
rect 4304 5324 4353 5352
rect 4304 5312 4310 5324
rect 4341 5321 4353 5324
rect 4387 5321 4399 5355
rect 4341 5315 4399 5321
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2363 5188 2605 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5185 3939 5219
rect 4356 5216 4384 5315
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 7006 5352 7012 5364
rect 6595 5324 7012 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7098 5312 7104 5364
rect 7156 5312 7162 5364
rect 9306 5312 9312 5364
rect 9364 5312 9370 5364
rect 5276 5256 5764 5284
rect 5276 5225 5304 5256
rect 5736 5228 5764 5256
rect 6822 5244 6828 5296
rect 6880 5284 6886 5296
rect 6880 5256 6960 5284
rect 6880 5244 6886 5256
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4356 5188 4721 5216
rect 3881 5179 3939 5185
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1673 5151 1731 5157
rect 1673 5148 1685 5151
rect 1452 5120 1685 5148
rect 1452 5108 1458 5120
rect 1673 5117 1685 5120
rect 1719 5117 1731 5151
rect 3896 5148 3924 5179
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5368 5148 5396 5176
rect 3896 5120 5396 5148
rect 5460 5148 5488 5179
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 6932 5225 6960 5256
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7116 5216 7144 5312
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8174 5287 8232 5293
rect 8174 5284 8186 5287
rect 8076 5256 8186 5284
rect 8076 5244 8082 5256
rect 8174 5253 8186 5256
rect 8220 5253 8232 5287
rect 8174 5247 8232 5253
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 9401 5287 9459 5293
rect 9401 5284 9413 5287
rect 8536 5256 9413 5284
rect 8536 5244 8542 5256
rect 9401 5253 9413 5256
rect 9447 5253 9459 5287
rect 9401 5247 9459 5253
rect 9585 5287 9643 5293
rect 9585 5253 9597 5287
rect 9631 5284 9643 5287
rect 10042 5284 10048 5296
rect 9631 5256 10048 5284
rect 9631 5253 9643 5256
rect 9585 5247 9643 5253
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 7116 5188 7205 5216
rect 7009 5179 7067 5185
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7834 5216 7840 5228
rect 7515 5188 7840 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 5626 5148 5632 5160
rect 5460 5120 5632 5148
rect 1673 5111 1731 5117
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 7024 5148 7052 5179
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 7282 5148 7288 5160
rect 6135 5120 7288 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 7374 5108 7380 5160
rect 7432 5108 7438 5160
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 7101 5083 7159 5089
rect 5316 5052 6684 5080
rect 5316 5040 5322 5052
rect 2406 4972 2412 5024
rect 2464 4972 2470 5024
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3844 4984 3985 5012
rect 3844 4972 3850 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 3973 4975 4031 4981
rect 4893 5015 4951 5021
rect 4893 4981 4905 5015
rect 4939 5012 4951 5015
rect 5074 5012 5080 5024
rect 4939 4984 5080 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 5353 5015 5411 5021
rect 5353 5012 5365 5015
rect 5224 4984 5365 5012
rect 5224 4972 5230 4984
rect 5353 4981 5365 4984
rect 5399 4981 5411 5015
rect 5353 4975 5411 4981
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 6362 5012 6368 5024
rect 5500 4984 6368 5012
rect 5500 4972 5506 4984
rect 6362 4972 6368 4984
rect 6420 5012 6426 5024
rect 6546 5012 6552 5024
rect 6420 4984 6552 5012
rect 6420 4972 6426 4984
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 6656 5012 6684 5052
rect 7101 5049 7113 5083
rect 7147 5080 7159 5083
rect 7576 5080 7604 5111
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 7147 5052 7604 5080
rect 7147 5049 7159 5052
rect 7101 5043 7159 5049
rect 7116 5012 7144 5043
rect 6656 4984 7144 5012
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 8294 5012 8300 5024
rect 7883 4984 8300 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 1104 4922 10028 4944
rect 1104 4870 2065 4922
rect 2117 4870 2129 4922
rect 2181 4870 2193 4922
rect 2245 4870 2257 4922
rect 2309 4870 2321 4922
rect 2373 4870 4296 4922
rect 4348 4870 4360 4922
rect 4412 4870 4424 4922
rect 4476 4870 4488 4922
rect 4540 4870 4552 4922
rect 4604 4870 6527 4922
rect 6579 4870 6591 4922
rect 6643 4870 6655 4922
rect 6707 4870 6719 4922
rect 6771 4870 6783 4922
rect 6835 4870 8758 4922
rect 8810 4870 8822 4922
rect 8874 4870 8886 4922
rect 8938 4870 8950 4922
rect 9002 4870 9014 4922
rect 9066 4870 10028 4922
rect 1104 4848 10028 4870
rect 1394 4768 1400 4820
rect 1452 4768 1458 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5902 4808 5908 4820
rect 5132 4780 5908 4808
rect 5132 4768 5138 4780
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 7024 4780 7420 4808
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 5994 4740 6000 4752
rect 4663 4712 6000 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5442 4672 5448 4684
rect 5316 4644 5448 4672
rect 5316 4632 5322 4644
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 7024 4681 7052 4780
rect 7392 4740 7420 4780
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7708 4780 7849 4808
rect 7708 4768 7714 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 7837 4771 7895 4777
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 9048 4740 9076 4771
rect 7392 4712 9076 4740
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3878 4604 3884 4616
rect 2823 4576 3884 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4798 4604 4804 4616
rect 4755 4576 4804 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 1946 4496 1952 4548
rect 2004 4536 2010 4548
rect 2510 4539 2568 4545
rect 2510 4536 2522 4539
rect 2004 4508 2522 4536
rect 2004 4496 2010 4508
rect 2510 4505 2522 4508
rect 2556 4505 2568 4539
rect 2510 4499 2568 4505
rect 4430 4496 4436 4548
rect 4488 4536 4494 4548
rect 4724 4536 4752 4567
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4604 5043 4607
rect 5074 4604 5080 4616
rect 5031 4576 5080 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5276 4545 5304 4632
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 5399 4576 5488 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 4488 4508 4752 4536
rect 5261 4539 5319 4545
rect 4488 4496 4494 4508
rect 5261 4505 5273 4539
rect 5307 4505 5319 4539
rect 5261 4499 5319 4505
rect 5460 4480 5488 4576
rect 6288 4576 7205 4604
rect 6288 4548 6316 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7340 4576 7665 4604
rect 7340 4564 7346 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 7653 4567 7711 4573
rect 8404 4576 9597 4604
rect 6270 4496 6276 4548
rect 6328 4496 6334 4548
rect 7006 4496 7012 4548
rect 7064 4496 7070 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 8404 4545 8432 4576
rect 9585 4573 9597 4576
rect 9631 4604 9643 4607
rect 9766 4604 9772 4616
rect 9631 4576 9772 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7156 4508 7481 4536
rect 7156 4496 7162 4508
rect 7469 4505 7481 4508
rect 7515 4505 7527 4539
rect 7469 4499 7527 4505
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4505 8447 4539
rect 8389 4499 8447 4505
rect 8757 4539 8815 4545
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 8803 4508 9904 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 4798 4428 4804 4480
rect 4856 4468 4862 4480
rect 5077 4471 5135 4477
rect 5077 4468 5089 4471
rect 4856 4440 5089 4468
rect 4856 4428 4862 4440
rect 5077 4437 5089 4440
rect 5123 4437 5135 4471
rect 5077 4431 5135 4437
rect 5442 4428 5448 4480
rect 5500 4428 5506 4480
rect 7024 4468 7052 4496
rect 8404 4468 8432 4499
rect 9876 4480 9904 4508
rect 7024 4440 8432 4468
rect 9858 4428 9864 4480
rect 9916 4428 9922 4480
rect 1104 4378 10028 4400
rect 1104 4326 2725 4378
rect 2777 4326 2789 4378
rect 2841 4326 2853 4378
rect 2905 4326 2917 4378
rect 2969 4326 2981 4378
rect 3033 4326 4956 4378
rect 5008 4326 5020 4378
rect 5072 4326 5084 4378
rect 5136 4326 5148 4378
rect 5200 4326 5212 4378
rect 5264 4326 7187 4378
rect 7239 4326 7251 4378
rect 7303 4326 7315 4378
rect 7367 4326 7379 4378
rect 7431 4326 7443 4378
rect 7495 4326 9418 4378
rect 9470 4326 9482 4378
rect 9534 4326 9546 4378
rect 9598 4326 9610 4378
rect 9662 4326 9674 4378
rect 9726 4326 10028 4378
rect 1104 4304 10028 4326
rect 2406 4264 2412 4276
rect 1780 4236 2412 4264
rect 1780 4137 1808 4236
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 4430 4224 4436 4276
rect 4488 4224 4494 4276
rect 4709 4267 4767 4273
rect 4709 4233 4721 4267
rect 4755 4233 4767 4267
rect 4709 4227 4767 4233
rect 2225 4199 2283 4205
rect 2225 4165 2237 4199
rect 2271 4196 2283 4199
rect 2271 4168 2360 4196
rect 2271 4165 2283 4168
rect 2225 4159 2283 4165
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4097 1547 4131
rect 1489 4091 1547 4097
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4097 1823 4131
rect 1765 4091 1823 4097
rect 1504 4060 1532 4091
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1504 4032 2053 4060
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2332 4060 2360 4168
rect 2424 4168 4016 4196
rect 2424 4137 2452 4168
rect 3988 4140 4016 4168
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 3786 4128 3792 4140
rect 2731 4100 3792 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 4448 4128 4476 4224
rect 4387 4100 4476 4128
rect 4724 4128 4752 4227
rect 5350 4224 5356 4276
rect 5408 4224 5414 4276
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 6270 4264 6276 4276
rect 5960 4236 6276 4264
rect 5960 4224 5966 4236
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 7006 4264 7012 4276
rect 6420 4236 7012 4264
rect 6420 4224 6426 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 8294 4224 8300 4276
rect 8352 4224 8358 4276
rect 9677 4267 9735 4273
rect 9677 4233 9689 4267
rect 9723 4264 9735 4267
rect 9766 4264 9772 4276
rect 9723 4236 9772 4264
rect 9723 4233 9735 4236
rect 9677 4227 9735 4233
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 5552 4196 5580 4224
rect 5460 4168 5580 4196
rect 8312 4196 8340 4224
rect 8312 4168 8432 4196
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4724 4100 5181 4128
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 5169 4097 5181 4100
rect 5215 4128 5227 4131
rect 5350 4128 5356 4140
rect 5215 4100 5356 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5460 4137 5488 4168
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4097 5503 4131
rect 5445 4091 5503 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6052 4100 6929 4128
rect 6052 4088 6058 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 7098 4088 7104 4140
rect 7156 4088 7162 4140
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 7984 4100 8309 4128
rect 7984 4088 7990 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8404 4128 8432 4168
rect 8553 4131 8611 4137
rect 8553 4128 8565 4131
rect 8404 4100 8565 4128
rect 8297 4091 8355 4097
rect 8553 4097 8565 4100
rect 8599 4097 8611 4131
rect 8553 4091 8611 4097
rect 2869 4063 2927 4069
rect 2869 4060 2881 4063
rect 2332 4032 2881 4060
rect 2041 4023 2099 4029
rect 2869 4029 2881 4032
rect 2915 4029 2927 4063
rect 2869 4023 2927 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 3528 3936 3556 4023
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 4212 4032 4445 4060
rect 4212 4020 4218 4032
rect 4433 4029 4445 4032
rect 4479 4060 4491 4063
rect 4522 4060 4528 4072
rect 4479 4032 4528 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 6089 4063 6147 4069
rect 6089 4060 6101 4063
rect 4908 4032 6101 4060
rect 4908 3936 4936 4032
rect 6089 4029 6101 4032
rect 6135 4029 6147 4063
rect 6089 4023 6147 4029
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6328 4032 6837 4060
rect 6328 4020 6334 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 6362 3992 6368 4004
rect 5092 3964 6368 3992
rect 5092 3936 5120 3964
rect 6362 3952 6368 3964
rect 6420 3992 6426 4004
rect 7024 3992 7052 4023
rect 6420 3964 7052 3992
rect 6420 3952 6426 3964
rect 1670 3884 1676 3936
rect 1728 3884 1734 3936
rect 1946 3884 1952 3936
rect 2004 3884 2010 3936
rect 2498 3884 2504 3936
rect 2556 3884 2562 3936
rect 3510 3884 3516 3936
rect 3568 3884 3574 3936
rect 4890 3884 4896 3936
rect 4948 3884 4954 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5074 3924 5080 3936
rect 5031 3896 5080 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5316 3896 5549 3924
rect 5316 3884 5322 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 7282 3884 7288 3936
rect 7340 3884 7346 3936
rect 1104 3834 10028 3856
rect 1104 3782 2065 3834
rect 2117 3782 2129 3834
rect 2181 3782 2193 3834
rect 2245 3782 2257 3834
rect 2309 3782 2321 3834
rect 2373 3782 4296 3834
rect 4348 3782 4360 3834
rect 4412 3782 4424 3834
rect 4476 3782 4488 3834
rect 4540 3782 4552 3834
rect 4604 3782 6527 3834
rect 6579 3782 6591 3834
rect 6643 3782 6655 3834
rect 6707 3782 6719 3834
rect 6771 3782 6783 3834
rect 6835 3782 8758 3834
rect 8810 3782 8822 3834
rect 8874 3782 8886 3834
rect 8938 3782 8950 3834
rect 9002 3782 9014 3834
rect 9066 3782 10028 3834
rect 1104 3760 10028 3782
rect 4065 3723 4123 3729
rect 2148 3692 3924 3720
rect 1578 3544 1584 3596
rect 1636 3584 1642 3596
rect 2148 3593 2176 3692
rect 3786 3612 3792 3664
rect 3844 3612 3850 3664
rect 3896 3596 3924 3692
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 4154 3720 4160 3732
rect 4111 3692 4160 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 4948 3692 7021 3720
rect 4948 3680 4954 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 7009 3683 7067 3689
rect 7282 3680 7288 3732
rect 7340 3680 7346 3732
rect 5534 3612 5540 3664
rect 5592 3612 5598 3664
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1636 3556 2145 3584
rect 1636 3544 1642 3556
rect 2133 3553 2145 3556
rect 2179 3553 2191 3587
rect 2133 3547 2191 3553
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 7300 3584 7328 3680
rect 3936 3556 5672 3584
rect 7300 3556 7420 3584
rect 3936 3544 3942 3556
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2389 3519 2447 3525
rect 2389 3516 2401 3519
rect 1728 3488 2401 3516
rect 1728 3476 1734 3488
rect 2389 3485 2401 3488
rect 2435 3485 2447 3519
rect 2389 3479 2447 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 1765 3451 1823 3457
rect 1765 3417 1777 3451
rect 1811 3448 1823 3451
rect 3988 3448 4016 3479
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4244 3519 4302 3525
rect 4244 3516 4256 3519
rect 4120 3488 4256 3516
rect 4120 3476 4126 3488
rect 4244 3485 4256 3488
rect 4290 3485 4302 3519
rect 4244 3479 4302 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4561 3519 4619 3525
rect 4561 3516 4573 3519
rect 4433 3479 4491 3485
rect 4540 3485 4573 3516
rect 4607 3485 4619 3519
rect 4540 3479 4619 3485
rect 4154 3448 4160 3460
rect 1811 3420 2774 3448
rect 3988 3420 4160 3448
rect 1811 3417 1823 3420
rect 1765 3411 1823 3417
rect 1486 3340 1492 3392
rect 1544 3340 1550 3392
rect 2746 3380 2774 3420
rect 4154 3408 4160 3420
rect 4212 3408 4218 3460
rect 4341 3451 4399 3457
rect 4341 3417 4353 3451
rect 4387 3417 4399 3451
rect 4341 3411 4399 3417
rect 3510 3380 3516 3392
rect 2746 3352 3516 3380
rect 3510 3340 3516 3352
rect 3568 3380 3574 3392
rect 4356 3380 4384 3411
rect 4448 3392 4476 3479
rect 4540 3448 4568 3479
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4985 3519 5043 3525
rect 4985 3516 4997 3519
rect 4856 3488 4997 3516
rect 4856 3476 4862 3488
rect 4985 3485 4997 3488
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 5132 3488 5181 3516
rect 5132 3476 5138 3488
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5258 3476 5264 3528
rect 5316 3476 5322 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5399 3488 5488 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 4890 3448 4896 3460
rect 4540 3420 4896 3448
rect 4540 3392 4568 3420
rect 4890 3408 4896 3420
rect 4948 3408 4954 3460
rect 3568 3352 4384 3380
rect 3568 3340 3574 3352
rect 4430 3340 4436 3392
rect 4488 3340 4494 3392
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 5460 3380 5488 3488
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 5644 3525 5672 3556
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 5718 3516 5724 3528
rect 5675 3488 5724 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6270 3476 6276 3528
rect 6328 3476 6334 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7392 3525 7420 3556
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 6972 3488 7297 3516
rect 6972 3476 6978 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 7791 3488 8953 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9088 3488 9505 3516
rect 9088 3476 9094 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 5552 3448 5580 3476
rect 5874 3451 5932 3457
rect 5874 3448 5886 3451
rect 5552 3420 5886 3448
rect 5874 3417 5886 3420
rect 5920 3417 5932 3451
rect 5874 3411 5932 3417
rect 6288 3448 6316 3476
rect 7653 3451 7711 3457
rect 7653 3448 7665 3451
rect 6288 3420 7665 3448
rect 6288 3380 6316 3420
rect 7653 3417 7665 3420
rect 7699 3417 7711 3451
rect 7653 3411 7711 3417
rect 8389 3451 8447 3457
rect 8389 3417 8401 3451
rect 8435 3448 8447 3451
rect 8570 3448 8576 3460
rect 8435 3420 8576 3448
rect 8435 3417 8447 3420
rect 8389 3411 8447 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 5460 3352 6316 3380
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 7558 3380 7564 3392
rect 7147 3352 7564 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 1104 3290 10028 3312
rect 1104 3238 2725 3290
rect 2777 3238 2789 3290
rect 2841 3238 2853 3290
rect 2905 3238 2917 3290
rect 2969 3238 2981 3290
rect 3033 3238 4956 3290
rect 5008 3238 5020 3290
rect 5072 3238 5084 3290
rect 5136 3238 5148 3290
rect 5200 3238 5212 3290
rect 5264 3238 7187 3290
rect 7239 3238 7251 3290
rect 7303 3238 7315 3290
rect 7367 3238 7379 3290
rect 7431 3238 7443 3290
rect 7495 3238 9418 3290
rect 9470 3238 9482 3290
rect 9534 3238 9546 3290
rect 9598 3238 9610 3290
rect 9662 3238 9674 3290
rect 9726 3238 10028 3290
rect 1104 3216 10028 3238
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3878 3176 3884 3188
rect 3099 3148 3884 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4522 3176 4528 3188
rect 4264 3148 4528 3176
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 4264 3108 4292 3148
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 6818 3179 6876 3185
rect 6818 3145 6830 3179
rect 6864 3176 6876 3179
rect 6914 3176 6920 3188
rect 6864 3148 6920 3176
rect 6864 3145 6876 3148
rect 6818 3139 6876 3145
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 7834 3176 7840 3188
rect 7248 3148 7840 3176
rect 7248 3136 7254 3148
rect 7834 3136 7840 3148
rect 7892 3176 7898 3188
rect 7892 3148 8064 3176
rect 7892 3136 7898 3148
rect 1811 3080 4292 3108
rect 4341 3111 4399 3117
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4614 3108 4620 3120
rect 4387 3080 4620 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4614 3068 4620 3080
rect 4672 3068 4678 3120
rect 5460 3080 5672 3108
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2409 3043 2467 3049
rect 2409 3009 2421 3043
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 2056 2972 2084 3003
rect 1360 2944 2084 2972
rect 2424 2972 2452 3003
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5460 3040 5488 3080
rect 4488 3012 5488 3040
rect 4488 3000 4494 3012
rect 5534 3000 5540 3052
rect 5592 3049 5598 3052
rect 5592 3003 5604 3049
rect 5644 3040 5672 3080
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 8036 3108 8064 3148
rect 8941 3111 8999 3117
rect 8941 3108 8953 3111
rect 5776 3080 7972 3108
rect 8036 3080 8953 3108
rect 5776 3068 5782 3080
rect 5828 3049 5856 3080
rect 5813 3043 5871 3049
rect 5644 3012 5764 3040
rect 5592 3000 5598 3003
rect 5736 2972 5764 3012
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6089 3043 6147 3049
rect 6089 3009 6101 3043
rect 6135 3040 6147 3043
rect 6270 3040 6276 3052
rect 6135 3012 6276 3040
rect 6135 3009 6147 3012
rect 6089 3003 6147 3009
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6420 3012 6653 3040
rect 6420 3000 6426 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 6012 2972 6040 3000
rect 6748 2972 6776 3003
rect 2424 2944 2774 2972
rect 5736 2944 5856 2972
rect 6012 2944 6776 2972
rect 6932 2972 6960 3003
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 7098 3000 7104 3052
rect 7156 3000 7162 3052
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7300 3049 7328 3080
rect 7944 3052 7972 3080
rect 8941 3077 8953 3080
rect 8987 3077 8999 3111
rect 8941 3071 8999 3077
rect 7558 3049 7564 3052
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7552 3040 7564 3049
rect 7519 3012 7564 3040
rect 7285 3003 7343 3009
rect 7552 3003 7564 3012
rect 7558 3000 7564 3003
rect 7616 3000 7622 3052
rect 7926 3000 7932 3052
rect 7984 3000 7990 3052
rect 7116 2972 7144 3000
rect 6932 2944 7144 2972
rect 1360 2932 1366 2944
rect 2746 2904 2774 2944
rect 5828 2904 5856 2944
rect 5997 2907 6055 2913
rect 5997 2904 6009 2907
rect 2746 2876 4936 2904
rect 5828 2876 6009 2904
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 72 2808 1501 2836
rect 72 2796 78 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 1489 2799 1547 2805
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4433 2839 4491 2845
rect 4433 2836 4445 2839
rect 4304 2808 4445 2836
rect 4304 2796 4310 2808
rect 4433 2805 4445 2808
rect 4479 2836 4491 2839
rect 4706 2836 4712 2848
rect 4479 2808 4712 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 4908 2836 4936 2876
rect 5997 2873 6009 2876
rect 6043 2904 6055 2907
rect 7208 2904 7236 3000
rect 6043 2876 7236 2904
rect 6043 2873 6055 2876
rect 5997 2867 6055 2873
rect 5626 2836 5632 2848
rect 4908 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 7190 2796 7196 2848
rect 7248 2796 7254 2848
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8260 2808 8677 2836
rect 8260 2796 8266 2808
rect 8665 2805 8677 2808
rect 8711 2836 8723 2839
rect 9030 2836 9036 2848
rect 8711 2808 9036 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9766 2836 9772 2848
rect 9263 2808 9772 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 1104 2746 10028 2768
rect 1104 2694 2065 2746
rect 2117 2694 2129 2746
rect 2181 2694 2193 2746
rect 2245 2694 2257 2746
rect 2309 2694 2321 2746
rect 2373 2694 4296 2746
rect 4348 2694 4360 2746
rect 4412 2694 4424 2746
rect 4476 2694 4488 2746
rect 4540 2694 4552 2746
rect 4604 2694 6527 2746
rect 6579 2694 6591 2746
rect 6643 2694 6655 2746
rect 6707 2694 6719 2746
rect 6771 2694 6783 2746
rect 6835 2694 8758 2746
rect 8810 2694 8822 2746
rect 8874 2694 8886 2746
rect 8938 2694 8950 2746
rect 9002 2694 9014 2746
rect 9066 2694 10028 2746
rect 1104 2672 10028 2694
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 4212 2604 4445 2632
rect 4212 2592 4218 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 6733 2499 6791 2505
rect 6733 2496 6745 2499
rect 4120 2468 5212 2496
rect 4120 2456 4126 2468
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2428 1547 2431
rect 1578 2428 1584 2440
rect 1535 2400 1584 2428
rect 1535 2397 1547 2400
rect 1489 2391 1547 2397
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1756 2431 1814 2437
rect 1756 2397 1768 2431
rect 1802 2428 1814 2431
rect 2498 2428 2504 2440
rect 1802 2400 2504 2428
rect 1802 2397 1814 2400
rect 1756 2391 1814 2397
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 2774 2320 2780 2372
rect 2832 2360 2838 2372
rect 3145 2363 3203 2369
rect 3145 2360 3157 2363
rect 2832 2332 3157 2360
rect 2832 2320 2838 2332
rect 3145 2329 3157 2332
rect 3191 2329 3203 2363
rect 3145 2323 3203 2329
rect 3513 2363 3571 2369
rect 3513 2329 3525 2363
rect 3559 2360 3571 2363
rect 3804 2360 3832 2391
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5184 2437 5212 2468
rect 5368 2468 6745 2496
rect 5368 2437 5396 2468
rect 6733 2465 6745 2468
rect 6779 2465 6791 2499
rect 6733 2459 6791 2465
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2496 7711 2499
rect 10962 2496 10968 2508
rect 7699 2468 10968 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 5169 2431 5227 2437
rect 4764 2400 5120 2428
rect 4764 2388 4770 2400
rect 3559 2332 3832 2360
rect 3559 2329 3571 2332
rect 3513 2323 3571 2329
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 3528 2292 3556 2323
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 4580 2332 4813 2360
rect 4580 2320 4586 2332
rect 4801 2329 4813 2332
rect 4847 2329 4859 2363
rect 5092 2360 5120 2400
rect 5169 2397 5181 2431
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 5684 2400 6377 2428
rect 5684 2388 5690 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7248 2400 7941 2428
rect 7248 2388 7254 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5092 2332 6101 2360
rect 4801 2323 4859 2329
rect 6089 2329 6101 2332
rect 6135 2360 6147 2363
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6135 2332 6561 2360
rect 6135 2329 6147 2332
rect 6089 2323 6147 2329
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6549 2323 6607 2329
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 8202 2360 8208 2372
rect 7423 2332 8208 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 2915 2264 3556 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 5810 2252 5816 2304
rect 5868 2252 5874 2304
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 7392 2292 7420 2323
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 6236 2264 7420 2292
rect 6236 2252 6242 2264
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 9030 2252 9036 2304
rect 9088 2252 9094 2304
rect 1104 2202 10028 2224
rect 1104 2150 2725 2202
rect 2777 2150 2789 2202
rect 2841 2150 2853 2202
rect 2905 2150 2917 2202
rect 2969 2150 2981 2202
rect 3033 2150 4956 2202
rect 5008 2150 5020 2202
rect 5072 2150 5084 2202
rect 5136 2150 5148 2202
rect 5200 2150 5212 2202
rect 5264 2150 7187 2202
rect 7239 2150 7251 2202
rect 7303 2150 7315 2202
rect 7367 2150 7379 2202
rect 7431 2150 7443 2202
rect 7495 2150 9418 2202
rect 9470 2150 9482 2202
rect 9534 2150 9546 2202
rect 9598 2150 9610 2202
rect 9662 2150 9674 2202
rect 9726 2150 10028 2202
rect 1104 2128 10028 2150
<< via1 >>
rect 2725 10854 2777 10906
rect 2789 10854 2841 10906
rect 2853 10854 2905 10906
rect 2917 10854 2969 10906
rect 2981 10854 3033 10906
rect 4956 10854 5008 10906
rect 5020 10854 5072 10906
rect 5084 10854 5136 10906
rect 5148 10854 5200 10906
rect 5212 10854 5264 10906
rect 7187 10854 7239 10906
rect 7251 10854 7303 10906
rect 7315 10854 7367 10906
rect 7379 10854 7431 10906
rect 7443 10854 7495 10906
rect 9418 10854 9470 10906
rect 9482 10854 9534 10906
rect 9546 10854 9598 10906
rect 9610 10854 9662 10906
rect 9674 10854 9726 10906
rect 2596 10752 2648 10804
rect 3056 10752 3108 10804
rect 3884 10752 3936 10804
rect 5816 10752 5868 10804
rect 7104 10752 7156 10804
rect 9312 10795 9364 10804
rect 9312 10761 9321 10795
rect 9321 10761 9355 10795
rect 9355 10761 9364 10795
rect 9312 10752 9364 10761
rect 2964 10616 3016 10668
rect 2596 10548 2648 10600
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4804 10616 4856 10668
rect 7656 10616 7708 10668
rect 8392 10548 8444 10600
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 3056 10412 3108 10464
rect 3240 10455 3292 10464
rect 3240 10421 3249 10455
rect 3249 10421 3283 10455
rect 3283 10421 3292 10455
rect 3240 10412 3292 10421
rect 7012 10412 7064 10464
rect 2065 10310 2117 10362
rect 2129 10310 2181 10362
rect 2193 10310 2245 10362
rect 2257 10310 2309 10362
rect 2321 10310 2373 10362
rect 4296 10310 4348 10362
rect 4360 10310 4412 10362
rect 4424 10310 4476 10362
rect 4488 10310 4540 10362
rect 4552 10310 4604 10362
rect 6527 10310 6579 10362
rect 6591 10310 6643 10362
rect 6655 10310 6707 10362
rect 6719 10310 6771 10362
rect 6783 10310 6835 10362
rect 8758 10310 8810 10362
rect 8822 10310 8874 10362
rect 8886 10310 8938 10362
rect 8950 10310 9002 10362
rect 9014 10310 9066 10362
rect 1308 10208 1360 10260
rect 3424 10208 3476 10260
rect 10324 10208 10376 10260
rect 3056 10183 3108 10192
rect 3056 10149 3065 10183
rect 3065 10149 3099 10183
rect 3099 10149 3108 10183
rect 3056 10140 3108 10149
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2504 10004 2556 10056
rect 4712 10004 4764 10056
rect 5356 10004 5408 10056
rect 5448 10047 5500 10056
rect 5448 10013 5457 10047
rect 5457 10013 5491 10047
rect 5491 10013 5500 10047
rect 5448 10004 5500 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 2228 9936 2280 9988
rect 5816 9936 5868 9988
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 7932 9936 7984 9988
rect 9772 9936 9824 9988
rect 4620 9868 4672 9920
rect 5540 9868 5592 9920
rect 5632 9868 5684 9920
rect 7012 9868 7064 9920
rect 7104 9868 7156 9920
rect 8024 9868 8076 9920
rect 8392 9868 8444 9920
rect 8944 9911 8996 9920
rect 8944 9877 8953 9911
rect 8953 9877 8987 9911
rect 8987 9877 8996 9911
rect 8944 9868 8996 9877
rect 2725 9766 2777 9818
rect 2789 9766 2841 9818
rect 2853 9766 2905 9818
rect 2917 9766 2969 9818
rect 2981 9766 3033 9818
rect 4956 9766 5008 9818
rect 5020 9766 5072 9818
rect 5084 9766 5136 9818
rect 5148 9766 5200 9818
rect 5212 9766 5264 9818
rect 7187 9766 7239 9818
rect 7251 9766 7303 9818
rect 7315 9766 7367 9818
rect 7379 9766 7431 9818
rect 7443 9766 7495 9818
rect 9418 9766 9470 9818
rect 9482 9766 9534 9818
rect 9546 9766 9598 9818
rect 9610 9766 9662 9818
rect 9674 9766 9726 9818
rect 1400 9664 1452 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 2228 9707 2280 9716
rect 2228 9673 2237 9707
rect 2237 9673 2271 9707
rect 2271 9673 2280 9707
rect 2228 9664 2280 9673
rect 4068 9664 4120 9716
rect 5540 9664 5592 9716
rect 5632 9664 5684 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 3240 9528 3292 9580
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3240 9392 3292 9444
rect 4620 9528 4672 9580
rect 4804 9528 4856 9580
rect 8392 9596 8444 9648
rect 8944 9596 8996 9648
rect 7104 9528 7156 9580
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7656 9460 7708 9512
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 9772 9392 9824 9444
rect 1768 9324 1820 9376
rect 2688 9324 2740 9376
rect 4068 9324 4120 9376
rect 4160 9324 4212 9376
rect 4712 9324 4764 9376
rect 6920 9324 6972 9376
rect 7104 9367 7156 9376
rect 7104 9333 7113 9367
rect 7113 9333 7147 9367
rect 7147 9333 7156 9367
rect 7104 9324 7156 9333
rect 8208 9324 8260 9376
rect 2065 9222 2117 9274
rect 2129 9222 2181 9274
rect 2193 9222 2245 9274
rect 2257 9222 2309 9274
rect 2321 9222 2373 9274
rect 4296 9222 4348 9274
rect 4360 9222 4412 9274
rect 4424 9222 4476 9274
rect 4488 9222 4540 9274
rect 4552 9222 4604 9274
rect 6527 9222 6579 9274
rect 6591 9222 6643 9274
rect 6655 9222 6707 9274
rect 6719 9222 6771 9274
rect 6783 9222 6835 9274
rect 8758 9222 8810 9274
rect 8822 9222 8874 9274
rect 8886 9222 8938 9274
rect 8950 9222 9002 9274
rect 9014 9222 9066 9274
rect 3056 9120 3108 9172
rect 4068 9120 4120 9172
rect 3240 9052 3292 9104
rect 5356 9052 5408 9104
rect 7840 9120 7892 9172
rect 7932 9163 7984 9172
rect 7932 9129 7941 9163
rect 7941 9129 7975 9163
rect 7975 9129 7984 9163
rect 7932 9120 7984 9129
rect 8116 9120 8168 9172
rect 2504 8984 2556 9036
rect 3792 8984 3844 9036
rect 4620 8984 4672 9036
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 4804 8916 4856 8968
rect 5448 8916 5500 8968
rect 8300 8984 8352 9036
rect 6092 8891 6144 8900
rect 6092 8857 6101 8891
rect 6101 8857 6135 8891
rect 6135 8857 6144 8891
rect 6092 8848 6144 8857
rect 2228 8780 2280 8832
rect 2688 8780 2740 8832
rect 4068 8780 4120 8832
rect 8024 8916 8076 8968
rect 8576 8984 8628 9036
rect 9772 8984 9824 9036
rect 7932 8848 7984 8900
rect 8484 8780 8536 8832
rect 9680 8848 9732 8900
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 2725 8678 2777 8730
rect 2789 8678 2841 8730
rect 2853 8678 2905 8730
rect 2917 8678 2969 8730
rect 2981 8678 3033 8730
rect 4956 8678 5008 8730
rect 5020 8678 5072 8730
rect 5084 8678 5136 8730
rect 5148 8678 5200 8730
rect 5212 8678 5264 8730
rect 7187 8678 7239 8730
rect 7251 8678 7303 8730
rect 7315 8678 7367 8730
rect 7379 8678 7431 8730
rect 7443 8678 7495 8730
rect 9418 8678 9470 8730
rect 9482 8678 9534 8730
rect 9546 8678 9598 8730
rect 9610 8678 9662 8730
rect 9674 8678 9726 8730
rect 1768 8576 1820 8628
rect 1860 8576 1912 8628
rect 2228 8576 2280 8628
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2504 8576 2556 8628
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 2504 8440 2556 8492
rect 3056 8576 3108 8628
rect 4804 8576 4856 8628
rect 5356 8576 5408 8628
rect 7840 8576 7892 8628
rect 9036 8576 9088 8628
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 3976 8508 4028 8560
rect 4712 8551 4764 8560
rect 4712 8517 4721 8551
rect 4721 8517 4755 8551
rect 4755 8517 4764 8551
rect 4712 8508 4764 8517
rect 5080 8483 5132 8492
rect 5080 8449 5114 8483
rect 5114 8449 5132 8483
rect 5080 8440 5132 8449
rect 9312 8440 9364 8492
rect 3332 8372 3384 8424
rect 9128 8372 9180 8424
rect 7932 8236 7984 8288
rect 2065 8134 2117 8186
rect 2129 8134 2181 8186
rect 2193 8134 2245 8186
rect 2257 8134 2309 8186
rect 2321 8134 2373 8186
rect 4296 8134 4348 8186
rect 4360 8134 4412 8186
rect 4424 8134 4476 8186
rect 4488 8134 4540 8186
rect 4552 8134 4604 8186
rect 6527 8134 6579 8186
rect 6591 8134 6643 8186
rect 6655 8134 6707 8186
rect 6719 8134 6771 8186
rect 6783 8134 6835 8186
rect 8758 8134 8810 8186
rect 8822 8134 8874 8186
rect 8886 8134 8938 8186
rect 8950 8134 9002 8186
rect 9014 8134 9066 8186
rect 940 8032 992 8084
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 3976 8032 4028 8084
rect 5080 8032 5132 8084
rect 6092 8032 6144 8084
rect 2412 7896 2464 7948
rect 2596 7828 2648 7880
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 3516 7828 3568 7880
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5908 7828 5960 7880
rect 7748 7964 7800 8016
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 7196 7896 7248 7948
rect 6368 7828 6420 7880
rect 6828 7828 6880 7880
rect 4068 7760 4120 7812
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 2412 7692 2464 7744
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 3424 7692 3476 7744
rect 6092 7692 6144 7744
rect 6276 7692 6328 7744
rect 7012 7692 7064 7744
rect 8392 7692 8444 7744
rect 9956 7692 10008 7744
rect 2725 7590 2777 7642
rect 2789 7590 2841 7642
rect 2853 7590 2905 7642
rect 2917 7590 2969 7642
rect 2981 7590 3033 7642
rect 4956 7590 5008 7642
rect 5020 7590 5072 7642
rect 5084 7590 5136 7642
rect 5148 7590 5200 7642
rect 5212 7590 5264 7642
rect 7187 7590 7239 7642
rect 7251 7590 7303 7642
rect 7315 7590 7367 7642
rect 7379 7590 7431 7642
rect 7443 7590 7495 7642
rect 9418 7590 9470 7642
rect 9482 7590 9534 7642
rect 9546 7590 9598 7642
rect 9610 7590 9662 7642
rect 9674 7590 9726 7642
rect 3056 7488 3108 7540
rect 3148 7488 3200 7540
rect 4804 7488 4856 7540
rect 7012 7488 7064 7540
rect 7932 7488 7984 7540
rect 8392 7488 8444 7540
rect 4620 7420 4672 7472
rect 5356 7420 5408 7472
rect 4160 7352 4212 7404
rect 4712 7327 4764 7336
rect 4712 7293 4721 7327
rect 4721 7293 4755 7327
rect 4755 7293 4764 7327
rect 4712 7284 4764 7293
rect 5448 7395 5500 7404
rect 5448 7361 5457 7395
rect 5457 7361 5491 7395
rect 5491 7361 5500 7395
rect 5448 7352 5500 7361
rect 6368 7352 6420 7404
rect 7472 7420 7524 7472
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 8024 7395 8076 7404
rect 7564 7327 7616 7336
rect 7564 7293 7573 7327
rect 7573 7293 7607 7327
rect 7607 7293 7616 7327
rect 7564 7284 7616 7293
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8392 7352 8444 7404
rect 6828 7216 6880 7268
rect 7656 7216 7708 7268
rect 4804 7148 4856 7200
rect 4988 7148 5040 7200
rect 7104 7191 7156 7200
rect 7104 7157 7113 7191
rect 7113 7157 7147 7191
rect 7147 7157 7156 7191
rect 7104 7148 7156 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 8208 7148 8260 7200
rect 2065 7046 2117 7098
rect 2129 7046 2181 7098
rect 2193 7046 2245 7098
rect 2257 7046 2309 7098
rect 2321 7046 2373 7098
rect 4296 7046 4348 7098
rect 4360 7046 4412 7098
rect 4424 7046 4476 7098
rect 4488 7046 4540 7098
rect 4552 7046 4604 7098
rect 6527 7046 6579 7098
rect 6591 7046 6643 7098
rect 6655 7046 6707 7098
rect 6719 7046 6771 7098
rect 6783 7046 6835 7098
rect 8758 7046 8810 7098
rect 8822 7046 8874 7098
rect 8886 7046 8938 7098
rect 8950 7046 9002 7098
rect 9014 7046 9066 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 3792 6944 3844 6996
rect 4252 6944 4304 6996
rect 4896 6944 4948 6996
rect 7104 6944 7156 6996
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 8024 6987 8076 6996
rect 8024 6953 8033 6987
rect 8033 6953 8067 6987
rect 8067 6953 8076 6987
rect 8024 6944 8076 6953
rect 8392 6944 8444 6996
rect 4620 6876 4672 6928
rect 1676 6740 1728 6792
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 940 6672 992 6724
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3332 6808 3384 6860
rect 4160 6808 4212 6860
rect 6920 6808 6972 6860
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 2504 6604 2556 6656
rect 3884 6604 3936 6656
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 4436 6740 4488 6792
rect 4988 6740 5040 6792
rect 6276 6740 6328 6792
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 8024 6808 8076 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 4160 6672 4212 6724
rect 7564 6672 7616 6724
rect 4528 6604 4580 6656
rect 5448 6604 5500 6656
rect 2725 6502 2777 6554
rect 2789 6502 2841 6554
rect 2853 6502 2905 6554
rect 2917 6502 2969 6554
rect 2981 6502 3033 6554
rect 4956 6502 5008 6554
rect 5020 6502 5072 6554
rect 5084 6502 5136 6554
rect 5148 6502 5200 6554
rect 5212 6502 5264 6554
rect 7187 6502 7239 6554
rect 7251 6502 7303 6554
rect 7315 6502 7367 6554
rect 7379 6502 7431 6554
rect 7443 6502 7495 6554
rect 9418 6502 9470 6554
rect 9482 6502 9534 6554
rect 9546 6502 9598 6554
rect 9610 6502 9662 6554
rect 9674 6502 9726 6554
rect 2044 6400 2096 6452
rect 2504 6400 2556 6452
rect 4344 6400 4396 6452
rect 4528 6443 4580 6452
rect 4528 6409 4537 6443
rect 4537 6409 4571 6443
rect 4571 6409 4580 6443
rect 4528 6400 4580 6409
rect 4712 6400 4764 6452
rect 6368 6400 6420 6452
rect 7012 6400 7064 6452
rect 7564 6400 7616 6452
rect 8116 6400 8168 6452
rect 8760 6400 8812 6452
rect 9312 6400 9364 6452
rect 3056 6332 3108 6384
rect 3608 6375 3660 6384
rect 3608 6341 3617 6375
rect 3617 6341 3651 6375
rect 3651 6341 3660 6375
rect 3608 6332 3660 6341
rect 3792 6332 3844 6384
rect 3516 6196 3568 6248
rect 3608 6196 3660 6248
rect 3884 6264 3936 6316
rect 4344 6264 4396 6316
rect 4528 6264 4580 6316
rect 4712 6264 4764 6316
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 5356 6264 5408 6316
rect 8208 6332 8260 6384
rect 4252 6196 4304 6248
rect 4436 6128 4488 6180
rect 4896 6196 4948 6248
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 5448 6196 5500 6205
rect 7840 6196 7892 6248
rect 7932 6196 7984 6248
rect 7012 6128 7064 6180
rect 3976 6060 4028 6112
rect 4344 6060 4396 6112
rect 4712 6060 4764 6112
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 5724 6103 5776 6112
rect 5724 6069 5733 6103
rect 5733 6069 5767 6103
rect 5767 6069 5776 6103
rect 5724 6060 5776 6069
rect 2065 5958 2117 6010
rect 2129 5958 2181 6010
rect 2193 5958 2245 6010
rect 2257 5958 2309 6010
rect 2321 5958 2373 6010
rect 4296 5958 4348 6010
rect 4360 5958 4412 6010
rect 4424 5958 4476 6010
rect 4488 5958 4540 6010
rect 4552 5958 4604 6010
rect 6527 5958 6579 6010
rect 6591 5958 6643 6010
rect 6655 5958 6707 6010
rect 6719 5958 6771 6010
rect 6783 5958 6835 6010
rect 8758 5958 8810 6010
rect 8822 5958 8874 6010
rect 8886 5958 8938 6010
rect 8950 5958 9002 6010
rect 9014 5958 9066 6010
rect 3424 5856 3476 5908
rect 3976 5856 4028 5908
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 7840 5856 7892 5908
rect 8024 5856 8076 5908
rect 9312 5788 9364 5840
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3884 5652 3936 5704
rect 1400 5584 1452 5636
rect 3516 5584 3568 5636
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 4988 5627 5040 5636
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 4160 5516 4212 5568
rect 4252 5559 4304 5568
rect 4252 5525 4277 5559
rect 4277 5525 4304 5559
rect 4252 5516 4304 5525
rect 4712 5516 4764 5568
rect 4988 5593 5013 5627
rect 5013 5593 5040 5627
rect 4988 5584 5040 5593
rect 5172 5516 5224 5568
rect 5356 5516 5408 5568
rect 5632 5516 5684 5568
rect 6552 5652 6604 5704
rect 7564 5652 7616 5704
rect 6828 5516 6880 5568
rect 7012 5516 7064 5568
rect 8024 5559 8076 5568
rect 8024 5525 8033 5559
rect 8033 5525 8067 5559
rect 8067 5525 8076 5559
rect 8024 5516 8076 5525
rect 2725 5414 2777 5466
rect 2789 5414 2841 5466
rect 2853 5414 2905 5466
rect 2917 5414 2969 5466
rect 2981 5414 3033 5466
rect 4956 5414 5008 5466
rect 5020 5414 5072 5466
rect 5084 5414 5136 5466
rect 5148 5414 5200 5466
rect 5212 5414 5264 5466
rect 7187 5414 7239 5466
rect 7251 5414 7303 5466
rect 7315 5414 7367 5466
rect 7379 5414 7431 5466
rect 7443 5414 7495 5466
rect 9418 5414 9470 5466
rect 9482 5414 9534 5466
rect 9546 5414 9598 5466
rect 9610 5414 9662 5466
rect 9674 5414 9726 5466
rect 4252 5312 4304 5364
rect 6276 5312 6328 5364
rect 7012 5312 7064 5364
rect 7104 5312 7156 5364
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 6828 5244 6880 5296
rect 1400 5108 1452 5160
rect 5356 5176 5408 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 8024 5244 8076 5296
rect 8484 5244 8536 5296
rect 10048 5244 10100 5296
rect 5632 5151 5684 5160
rect 5632 5117 5641 5151
rect 5641 5117 5675 5151
rect 5675 5117 5684 5151
rect 5632 5108 5684 5117
rect 7840 5176 7892 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 7288 5108 7340 5160
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 5264 5040 5316 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 3792 4972 3844 5024
rect 5080 4972 5132 5024
rect 5172 4972 5224 5024
rect 5448 4972 5500 5024
rect 6368 4972 6420 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 8300 4972 8352 5024
rect 2065 4870 2117 4922
rect 2129 4870 2181 4922
rect 2193 4870 2245 4922
rect 2257 4870 2309 4922
rect 2321 4870 2373 4922
rect 4296 4870 4348 4922
rect 4360 4870 4412 4922
rect 4424 4870 4476 4922
rect 4488 4870 4540 4922
rect 4552 4870 4604 4922
rect 6527 4870 6579 4922
rect 6591 4870 6643 4922
rect 6655 4870 6707 4922
rect 6719 4870 6771 4922
rect 6783 4870 6835 4922
rect 8758 4870 8810 4922
rect 8822 4870 8874 4922
rect 8886 4870 8938 4922
rect 8950 4870 9002 4922
rect 9014 4870 9066 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 5080 4768 5132 4820
rect 5908 4768 5960 4820
rect 6000 4700 6052 4752
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5264 4632 5316 4684
rect 5448 4632 5500 4684
rect 7656 4768 7708 4820
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 3884 4564 3936 4616
rect 4528 4607 4580 4616
rect 4528 4573 4537 4607
rect 4537 4573 4571 4607
rect 4571 4573 4580 4607
rect 4528 4564 4580 4573
rect 1952 4496 2004 4548
rect 4436 4496 4488 4548
rect 4804 4564 4856 4616
rect 5080 4564 5132 4616
rect 7288 4564 7340 4616
rect 6276 4496 6328 4548
rect 7012 4496 7064 4548
rect 7104 4496 7156 4548
rect 9772 4564 9824 4616
rect 4804 4428 4856 4480
rect 5448 4428 5500 4480
rect 9864 4428 9916 4480
rect 2725 4326 2777 4378
rect 2789 4326 2841 4378
rect 2853 4326 2905 4378
rect 2917 4326 2969 4378
rect 2981 4326 3033 4378
rect 4956 4326 5008 4378
rect 5020 4326 5072 4378
rect 5084 4326 5136 4378
rect 5148 4326 5200 4378
rect 5212 4326 5264 4378
rect 7187 4326 7239 4378
rect 7251 4326 7303 4378
rect 7315 4326 7367 4378
rect 7379 4326 7431 4378
rect 7443 4326 7495 4378
rect 9418 4326 9470 4378
rect 9482 4326 9534 4378
rect 9546 4326 9598 4378
rect 9610 4326 9662 4378
rect 9674 4326 9726 4378
rect 2412 4224 2464 4276
rect 4436 4224 4488 4276
rect 3792 4088 3844 4140
rect 3976 4088 4028 4140
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 5540 4224 5592 4276
rect 5908 4224 5960 4276
rect 6276 4224 6328 4276
rect 6368 4224 6420 4276
rect 7012 4224 7064 4276
rect 8300 4224 8352 4276
rect 9772 4224 9824 4276
rect 5356 4088 5408 4140
rect 6000 4088 6052 4140
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 7932 4088 7984 4140
rect 4160 4020 4212 4072
rect 4528 4020 4580 4072
rect 6276 4020 6328 4072
rect 6368 3952 6420 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 2504 3927 2556 3936
rect 2504 3893 2513 3927
rect 2513 3893 2547 3927
rect 2547 3893 2556 3927
rect 2504 3884 2556 3893
rect 3516 3884 3568 3936
rect 4896 3884 4948 3936
rect 5080 3884 5132 3936
rect 5264 3884 5316 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 2065 3782 2117 3834
rect 2129 3782 2181 3834
rect 2193 3782 2245 3834
rect 2257 3782 2309 3834
rect 2321 3782 2373 3834
rect 4296 3782 4348 3834
rect 4360 3782 4412 3834
rect 4424 3782 4476 3834
rect 4488 3782 4540 3834
rect 4552 3782 4604 3834
rect 6527 3782 6579 3834
rect 6591 3782 6643 3834
rect 6655 3782 6707 3834
rect 6719 3782 6771 3834
rect 6783 3782 6835 3834
rect 8758 3782 8810 3834
rect 8822 3782 8874 3834
rect 8886 3782 8938 3834
rect 8950 3782 9002 3834
rect 9014 3782 9066 3834
rect 1584 3544 1636 3596
rect 3792 3655 3844 3664
rect 3792 3621 3801 3655
rect 3801 3621 3835 3655
rect 3835 3621 3844 3655
rect 3792 3612 3844 3621
rect 4160 3680 4212 3732
rect 4896 3680 4948 3732
rect 7288 3680 7340 3732
rect 5540 3655 5592 3664
rect 5540 3621 5549 3655
rect 5549 3621 5583 3655
rect 5583 3621 5592 3655
rect 5540 3612 5592 3621
rect 3884 3544 3936 3596
rect 1676 3476 1728 3528
rect 4068 3476 4120 3528
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 4160 3408 4212 3460
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 4804 3476 4856 3528
rect 5080 3476 5132 3528
rect 5264 3519 5316 3528
rect 5264 3485 5273 3519
rect 5273 3485 5307 3519
rect 5307 3485 5316 3519
rect 5264 3476 5316 3485
rect 4896 3408 4948 3460
rect 3516 3340 3568 3349
rect 4436 3340 4488 3392
rect 4528 3340 4580 3392
rect 5540 3476 5592 3528
rect 5724 3476 5776 3528
rect 6276 3476 6328 3528
rect 6920 3476 6972 3528
rect 9036 3476 9088 3528
rect 8576 3408 8628 3460
rect 7564 3340 7616 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 2725 3238 2777 3290
rect 2789 3238 2841 3290
rect 2853 3238 2905 3290
rect 2917 3238 2969 3290
rect 2981 3238 3033 3290
rect 4956 3238 5008 3290
rect 5020 3238 5072 3290
rect 5084 3238 5136 3290
rect 5148 3238 5200 3290
rect 5212 3238 5264 3290
rect 7187 3238 7239 3290
rect 7251 3238 7303 3290
rect 7315 3238 7367 3290
rect 7379 3238 7431 3290
rect 7443 3238 7495 3290
rect 9418 3238 9470 3290
rect 9482 3238 9534 3290
rect 9546 3238 9598 3290
rect 9610 3238 9662 3290
rect 9674 3238 9726 3290
rect 3884 3136 3936 3188
rect 4528 3136 4580 3188
rect 6920 3136 6972 3188
rect 7196 3136 7248 3188
rect 7840 3136 7892 3188
rect 4620 3068 4672 3120
rect 1308 2932 1360 2984
rect 4436 3000 4488 3052
rect 5540 3043 5592 3052
rect 5540 3009 5558 3043
rect 5558 3009 5592 3043
rect 5540 3000 5592 3009
rect 5724 3068 5776 3120
rect 6000 3000 6052 3052
rect 6276 3000 6328 3052
rect 6368 3000 6420 3052
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7104 3000 7156 3052
rect 7196 3000 7248 3052
rect 7564 3043 7616 3052
rect 7564 3009 7598 3043
rect 7598 3009 7616 3043
rect 7564 3000 7616 3009
rect 7932 3000 7984 3052
rect 20 2796 72 2848
rect 4252 2796 4304 2848
rect 4712 2796 4764 2848
rect 5632 2796 5684 2848
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 8208 2796 8260 2848
rect 9036 2796 9088 2848
rect 9772 2796 9824 2848
rect 2065 2694 2117 2746
rect 2129 2694 2181 2746
rect 2193 2694 2245 2746
rect 2257 2694 2309 2746
rect 2321 2694 2373 2746
rect 4296 2694 4348 2746
rect 4360 2694 4412 2746
rect 4424 2694 4476 2746
rect 4488 2694 4540 2746
rect 4552 2694 4604 2746
rect 6527 2694 6579 2746
rect 6591 2694 6643 2746
rect 6655 2694 6707 2746
rect 6719 2694 6771 2746
rect 6783 2694 6835 2746
rect 8758 2694 8810 2746
rect 8822 2694 8874 2746
rect 8886 2694 8938 2746
rect 8950 2694 9002 2746
rect 9014 2694 9066 2746
rect 4160 2592 4212 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 4068 2456 4120 2508
rect 1584 2388 1636 2440
rect 2504 2388 2556 2440
rect 2780 2320 2832 2372
rect 4712 2388 4764 2440
rect 10968 2456 11020 2508
rect 4528 2320 4580 2372
rect 5632 2388 5684 2440
rect 7196 2388 7248 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 6184 2252 6236 2304
rect 8208 2320 8260 2372
rect 7748 2252 7800 2304
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9036 2252 9088 2261
rect 2725 2150 2777 2202
rect 2789 2150 2841 2202
rect 2853 2150 2905 2202
rect 2917 2150 2969 2202
rect 2981 2150 3033 2202
rect 4956 2150 5008 2202
rect 5020 2150 5072 2202
rect 5084 2150 5136 2202
rect 5148 2150 5200 2202
rect 5212 2150 5264 2202
rect 7187 2150 7239 2202
rect 7251 2150 7303 2202
rect 7315 2150 7367 2202
rect 7379 2150 7431 2202
rect 7443 2150 7495 2202
rect 9418 2150 9470 2202
rect 9482 2150 9534 2202
rect 9546 2150 9598 2202
rect 9610 2150 9662 2202
rect 9674 2150 9726 2202
<< metal2 >>
rect 1306 12534 1362 13334
rect 2594 12534 2650 13334
rect 3054 13016 3110 13025
rect 3054 12951 3110 12960
rect 1320 10266 1348 12534
rect 1582 11656 1638 11665
rect 1582 11591 1638 11600
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9722 1440 9998
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1504 9625 1532 10406
rect 1596 9654 1624 11591
rect 2608 10810 2636 12534
rect 2725 10908 3033 10917
rect 2725 10906 2731 10908
rect 2787 10906 2811 10908
rect 2867 10906 2891 10908
rect 2947 10906 2971 10908
rect 3027 10906 3033 10908
rect 2787 10854 2789 10906
rect 2969 10854 2971 10906
rect 2725 10852 2731 10854
rect 2787 10852 2811 10854
rect 2867 10852 2891 10854
rect 2947 10852 2971 10854
rect 3027 10852 3033 10854
rect 2725 10843 3033 10852
rect 3068 10810 3096 12951
rect 3882 12534 3938 13334
rect 5814 12534 5870 13334
rect 7102 12534 7158 13334
rect 9034 12534 9090 13334
rect 10322 12534 10378 13334
rect 3896 10810 3924 12534
rect 4956 10908 5264 10917
rect 4956 10906 4962 10908
rect 5018 10906 5042 10908
rect 5098 10906 5122 10908
rect 5178 10906 5202 10908
rect 5258 10906 5264 10908
rect 5018 10854 5020 10906
rect 5200 10854 5202 10906
rect 4956 10852 4962 10854
rect 5018 10852 5042 10854
rect 5098 10852 5122 10854
rect 5178 10852 5202 10854
rect 5258 10852 5264 10854
rect 4956 10843 5264 10852
rect 5828 10810 5856 12534
rect 7116 10810 7144 12534
rect 7187 10908 7495 10917
rect 7187 10906 7193 10908
rect 7249 10906 7273 10908
rect 7329 10906 7353 10908
rect 7409 10906 7433 10908
rect 7489 10906 7495 10908
rect 7249 10854 7251 10906
rect 7431 10854 7433 10906
rect 7187 10852 7193 10854
rect 7249 10852 7273 10854
rect 7329 10852 7353 10854
rect 7409 10852 7433 10854
rect 7489 10852 7495 10854
rect 7187 10843 7495 10852
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 8206 10704 8262 10713
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 7656 10668 7708 10674
rect 8206 10639 8262 10648
rect 7656 10610 7708 10616
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2065 10364 2373 10373
rect 2065 10362 2071 10364
rect 2127 10362 2151 10364
rect 2207 10362 2231 10364
rect 2287 10362 2311 10364
rect 2367 10362 2373 10364
rect 2127 10310 2129 10362
rect 2309 10310 2311 10362
rect 2065 10308 2071 10310
rect 2127 10308 2151 10310
rect 2207 10308 2231 10310
rect 2287 10308 2311 10310
rect 2367 10308 2373 10310
rect 2065 10299 2373 10308
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 9722 2268 9930
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 1584 9648 1636 9654
rect 1490 9616 1546 9625
rect 1584 9590 1636 9596
rect 1490 9551 1546 9560
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 8634 1808 9318
rect 2065 9276 2373 9285
rect 2065 9274 2071 9276
rect 2127 9274 2151 9276
rect 2207 9274 2231 9276
rect 2287 9274 2311 9276
rect 2367 9274 2373 9276
rect 2127 9222 2129 9274
rect 2309 9222 2311 9274
rect 2065 9220 2071 9222
rect 2127 9220 2151 9222
rect 2207 9220 2231 9222
rect 2287 9220 2311 9222
rect 2367 9220 2373 9222
rect 2065 9211 2373 9220
rect 2516 9042 2544 9998
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8634 1900 8842
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8634 2268 8774
rect 2516 8634 2544 8978
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 938 8256 994 8265
rect 938 8191 994 8200
rect 952 8090 980 8191
rect 940 8084 992 8090
rect 940 8026 992 8032
rect 1688 6798 1716 8366
rect 2065 8188 2373 8197
rect 2065 8186 2071 8188
rect 2127 8186 2151 8188
rect 2207 8186 2231 8188
rect 2287 8186 2311 8188
rect 2367 8186 2373 8188
rect 2127 8134 2129 8186
rect 2309 8134 2311 8186
rect 2065 8132 2071 8134
rect 2127 8132 2151 8134
rect 2207 8132 2231 8134
rect 2287 8132 2311 8134
rect 2367 8132 2373 8134
rect 2065 8123 2373 8132
rect 2424 7954 2452 8434
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2065 7100 2373 7109
rect 2065 7098 2071 7100
rect 2127 7098 2151 7100
rect 2207 7098 2231 7100
rect 2287 7098 2311 7100
rect 2367 7098 2373 7100
rect 2127 7046 2129 7098
rect 2309 7046 2311 7098
rect 2065 7044 2071 7046
rect 2127 7044 2151 7046
rect 2207 7044 2231 7046
rect 2287 7044 2311 7046
rect 2367 7044 2373 7046
rect 2065 7035 2373 7044
rect 2424 7002 2452 7686
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2516 6914 2544 8434
rect 2608 7886 2636 10542
rect 2976 10010 3004 10610
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3068 10198 3096 10406
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 2976 9982 3096 10010
rect 2725 9820 3033 9829
rect 2725 9818 2731 9820
rect 2787 9818 2811 9820
rect 2867 9818 2891 9820
rect 2947 9818 2971 9820
rect 3027 9818 3033 9820
rect 2787 9766 2789 9818
rect 2969 9766 2971 9818
rect 2725 9764 2731 9766
rect 2787 9764 2811 9766
rect 2867 9764 2891 9766
rect 2947 9764 2971 9766
rect 3027 9764 3033 9766
rect 2725 9755 3033 9764
rect 3068 9518 3096 9982
rect 3252 9586 3280 10406
rect 3436 10266 3464 10610
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 4080 9722 4108 10610
rect 4296 10364 4604 10373
rect 4296 10362 4302 10364
rect 4358 10362 4382 10364
rect 4438 10362 4462 10364
rect 4518 10362 4542 10364
rect 4598 10362 4604 10364
rect 4358 10310 4360 10362
rect 4540 10310 4542 10362
rect 4296 10308 4302 10310
rect 4358 10308 4382 10310
rect 4438 10308 4462 10310
rect 4518 10308 4542 10310
rect 4598 10308 4604 10310
rect 4296 10299 4604 10308
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4632 9586 4660 9862
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2700 8838 2728 9318
rect 3068 9178 3096 9454
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3252 9110 3280 9386
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4080 9178 4108 9318
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2725 8732 3033 8741
rect 2725 8730 2731 8732
rect 2787 8730 2811 8732
rect 2867 8730 2891 8732
rect 2947 8730 2971 8732
rect 3027 8730 3033 8732
rect 2787 8678 2789 8730
rect 2969 8678 2971 8730
rect 2725 8676 2731 8678
rect 2787 8676 2811 8678
rect 2867 8676 2891 8678
rect 2947 8676 2971 8678
rect 3027 8676 3033 8678
rect 2725 8667 3033 8676
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2725 7644 3033 7653
rect 2725 7642 2731 7644
rect 2787 7642 2811 7644
rect 2867 7642 2891 7644
rect 2947 7642 2971 7644
rect 3027 7642 3033 7644
rect 2787 7590 2789 7642
rect 2969 7590 2971 7642
rect 2725 7588 2731 7590
rect 2787 7588 2811 7590
rect 2867 7588 2891 7590
rect 2947 7588 2971 7590
rect 3027 7588 3033 7590
rect 2725 7579 3033 7588
rect 3068 7546 3096 8570
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3344 8090 3372 8366
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3516 7880 3568 7886
rect 3344 7840 3516 7868
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7546 3188 7686
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2516 6886 2728 6914
rect 1964 6854 2268 6882
rect 1964 6798 1992 6854
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6225 980 6666
rect 2056 6458 2084 6734
rect 2240 6662 2268 6854
rect 2700 6798 2728 6886
rect 3344 6866 3372 7840
rect 3516 7822 3568 7828
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3436 6798 3464 7686
rect 3804 7002 3832 8978
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3988 8090 4016 8502
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4080 7818 4108 8774
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4172 7698 4200 9318
rect 4296 9276 4604 9285
rect 4296 9274 4302 9276
rect 4358 9274 4382 9276
rect 4438 9274 4462 9276
rect 4518 9274 4542 9276
rect 4598 9274 4604 9276
rect 4358 9222 4360 9274
rect 4540 9222 4542 9274
rect 4296 9220 4302 9222
rect 4358 9220 4382 9222
rect 4438 9220 4462 9222
rect 4518 9220 4542 9222
rect 4598 9220 4604 9222
rect 4296 9211 4604 9220
rect 4632 9042 4660 9522
rect 4724 9382 4752 9998
rect 4816 9586 4844 10610
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6527 10364 6835 10373
rect 6527 10362 6533 10364
rect 6589 10362 6613 10364
rect 6669 10362 6693 10364
rect 6749 10362 6773 10364
rect 6829 10362 6835 10364
rect 6589 10310 6591 10362
rect 6771 10310 6773 10362
rect 6527 10308 6533 10310
rect 6589 10308 6613 10310
rect 6669 10308 6693 10310
rect 6749 10308 6773 10310
rect 6829 10308 6835 10310
rect 6527 10299 6835 10308
rect 7024 10062 7052 10406
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 4956 9820 5264 9829
rect 4956 9818 4962 9820
rect 5018 9818 5042 9820
rect 5098 9818 5122 9820
rect 5178 9818 5202 9820
rect 5258 9818 5264 9820
rect 5018 9766 5020 9818
rect 5200 9766 5202 9818
rect 4956 9764 4962 9766
rect 5018 9764 5042 9766
rect 5098 9764 5122 9766
rect 5178 9764 5202 9766
rect 5258 9764 5264 9766
rect 4956 9755 5264 9764
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4816 9058 4844 9522
rect 5368 9110 5396 9998
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4724 9030 4844 9058
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 4724 8566 4752 9030
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8634 4844 8910
rect 4956 8732 5264 8741
rect 4956 8730 4962 8732
rect 5018 8730 5042 8732
rect 5098 8730 5122 8732
rect 5178 8730 5202 8732
rect 5258 8730 5264 8732
rect 5018 8678 5020 8730
rect 5200 8678 5202 8730
rect 4956 8676 4962 8678
rect 5018 8676 5042 8678
rect 5098 8676 5122 8678
rect 5178 8676 5202 8678
rect 5258 8676 5264 8678
rect 4956 8667 5264 8676
rect 5368 8634 5396 9046
rect 5460 8974 5488 9998
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5552 9722 5580 9862
rect 5644 9722 5672 9862
rect 5828 9722 5856 9930
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 7024 9518 7052 9862
rect 7116 9586 7144 9862
rect 7187 9820 7495 9829
rect 7187 9818 7193 9820
rect 7249 9818 7273 9820
rect 7329 9818 7353 9820
rect 7409 9818 7433 9820
rect 7489 9818 7495 9820
rect 7249 9766 7251 9818
rect 7431 9766 7433 9818
rect 7187 9764 7193 9766
rect 7249 9764 7273 9766
rect 7329 9764 7353 9766
rect 7409 9764 7433 9766
rect 7489 9764 7495 9766
rect 7187 9755 7495 9764
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7668 9518 7696 10610
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6527 9276 6835 9285
rect 6527 9274 6533 9276
rect 6589 9274 6613 9276
rect 6669 9274 6693 9276
rect 6749 9274 6773 9276
rect 6829 9274 6835 9276
rect 6589 9222 6591 9274
rect 6771 9222 6773 9274
rect 6527 9220 6533 9222
rect 6589 9220 6613 9222
rect 6669 9220 6693 9222
rect 6749 9220 6773 9222
rect 6829 9220 6835 9222
rect 6527 9211 6835 9220
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4296 8188 4604 8197
rect 4296 8186 4302 8188
rect 4358 8186 4382 8188
rect 4438 8186 4462 8188
rect 4518 8186 4542 8188
rect 4598 8186 4604 8188
rect 4358 8134 4360 8186
rect 4540 8134 4542 8186
rect 4296 8132 4302 8134
rect 4358 8132 4382 8134
rect 4438 8132 4462 8134
rect 4518 8132 4542 8134
rect 4598 8132 4604 8134
rect 4296 8123 4604 8132
rect 4724 7954 4752 8502
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5092 8090 5120 8434
rect 6104 8090 6132 8842
rect 6527 8188 6835 8197
rect 6527 8186 6533 8188
rect 6589 8186 6613 8188
rect 6669 8186 6693 8188
rect 6749 8186 6773 8188
rect 6829 8186 6835 8188
rect 6589 8134 6591 8186
rect 6771 8134 6773 8186
rect 6527 8132 6533 8134
rect 6589 8132 6613 8134
rect 6669 8132 6693 8134
rect 6749 8132 6773 8134
rect 6829 8132 6835 8134
rect 6527 8123 6835 8132
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4080 7670 4200 7698
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3424 6792 3476 6798
rect 3476 6740 3556 6746
rect 3424 6734 3556 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6458 2544 6598
rect 2725 6556 3033 6565
rect 2725 6554 2731 6556
rect 2787 6554 2811 6556
rect 2867 6554 2891 6556
rect 2947 6554 2971 6556
rect 3027 6554 3033 6556
rect 2787 6502 2789 6554
rect 2969 6502 2971 6554
rect 2725 6500 2731 6502
rect 2787 6500 2811 6502
rect 2867 6500 2891 6502
rect 2947 6500 2971 6502
rect 3027 6500 3033 6502
rect 2725 6491 3033 6500
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 3068 6390 3096 6734
rect 3436 6718 3556 6734
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3528 6254 3556 6718
rect 3804 6390 3832 6938
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3608 6384 3660 6390
rect 3606 6352 3608 6361
rect 3792 6384 3844 6390
rect 3660 6352 3662 6361
rect 3792 6326 3844 6332
rect 3896 6322 3924 6598
rect 3606 6287 3662 6296
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3516 6248 3568 6254
rect 938 6216 994 6225
rect 3516 6190 3568 6196
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 938 6151 994 6160
rect 2065 6012 2373 6021
rect 2065 6010 2071 6012
rect 2127 6010 2151 6012
rect 2207 6010 2231 6012
rect 2287 6010 2311 6012
rect 2367 6010 2373 6012
rect 2127 5958 2129 6010
rect 2309 5958 2311 6010
rect 2065 5956 2071 5958
rect 2127 5956 2151 5958
rect 2207 5956 2231 5958
rect 2287 5956 2311 5958
rect 2367 5956 2373 5958
rect 2065 5947 2373 5956
rect 3528 5930 3556 6190
rect 3436 5914 3556 5930
rect 3424 5908 3556 5914
rect 3476 5902 3556 5908
rect 3424 5850 3476 5856
rect 3528 5642 3556 5902
rect 3620 5710 3648 6190
rect 3896 5794 3924 6258
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5914 4016 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5794 4108 7670
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4724 7426 4752 7890
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 4816 7546 4844 7822
rect 4956 7644 5264 7653
rect 4956 7642 4962 7644
rect 5018 7642 5042 7644
rect 5098 7642 5122 7644
rect 5178 7642 5202 7644
rect 5258 7642 5264 7644
rect 5018 7590 5020 7642
rect 5200 7590 5202 7642
rect 4956 7588 4962 7590
rect 5018 7588 5042 7590
rect 5098 7588 5122 7590
rect 5178 7588 5202 7590
rect 5258 7588 5264 7590
rect 4956 7579 5264 7588
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5356 7472 5408 7478
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 6866 4200 7346
rect 4296 7100 4604 7109
rect 4296 7098 4302 7100
rect 4358 7098 4382 7100
rect 4438 7098 4462 7100
rect 4518 7098 4542 7100
rect 4598 7098 4604 7100
rect 4358 7046 4360 7098
rect 4540 7046 4542 7098
rect 4296 7044 4302 7046
rect 4358 7044 4382 7046
rect 4438 7044 4462 7046
rect 4518 7044 4542 7046
rect 4598 7044 4604 7046
rect 4296 7035 4604 7044
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3804 5766 3924 5794
rect 3988 5766 4108 5794
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 1412 5166 1440 5578
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 1412 4826 1440 5102
rect 1872 5001 1900 5510
rect 2725 5468 3033 5477
rect 2725 5466 2731 5468
rect 2787 5466 2811 5468
rect 2867 5466 2891 5468
rect 2947 5466 2971 5468
rect 3027 5466 3033 5468
rect 2787 5414 2789 5466
rect 2969 5414 2971 5466
rect 2725 5412 2731 5414
rect 2787 5412 2811 5414
rect 2867 5412 2891 5414
rect 2947 5412 2971 5414
rect 3027 5412 3033 5414
rect 2725 5403 3033 5412
rect 3804 5030 3832 5766
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 2412 5024 2464 5030
rect 1858 4992 1914 5001
rect 2412 4966 2464 4972
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 1858 4927 1914 4936
rect 2065 4924 2373 4933
rect 2065 4922 2071 4924
rect 2127 4922 2151 4924
rect 2207 4922 2231 4924
rect 2287 4922 2311 4924
rect 2367 4922 2373 4924
rect 2127 4870 2129 4922
rect 2309 4870 2311 4922
rect 2065 4868 2071 4870
rect 2127 4868 2151 4870
rect 2207 4868 2231 4870
rect 2287 4868 2311 4870
rect 2367 4868 2373 4870
rect 2065 4859 2373 4868
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1964 3942 1992 4490
rect 2424 4282 2452 4966
rect 3896 4622 3924 5646
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 2725 4380 3033 4389
rect 2725 4378 2731 4380
rect 2787 4378 2811 4380
rect 2867 4378 2891 4380
rect 2947 4378 2971 4380
rect 3027 4378 3033 4380
rect 2787 4326 2789 4378
rect 2969 4326 2971 4378
rect 2725 4324 2731 4326
rect 2787 4324 2811 4326
rect 2867 4324 2891 4326
rect 2947 4324 2971 4326
rect 3027 4324 3033 4326
rect 2725 4315 3033 4324
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1320 800 1348 2926
rect 1504 1601 1532 3334
rect 1596 2446 1624 3538
rect 1688 3534 1716 3878
rect 2065 3836 2373 3845
rect 2065 3834 2071 3836
rect 2127 3834 2151 3836
rect 2207 3834 2231 3836
rect 2287 3834 2311 3836
rect 2367 3834 2373 3836
rect 2127 3782 2129 3834
rect 2309 3782 2311 3834
rect 2065 3780 2071 3782
rect 2127 3780 2151 3782
rect 2207 3780 2231 3782
rect 2287 3780 2311 3782
rect 2367 3780 2373 3782
rect 2065 3771 2373 3780
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2065 2748 2373 2757
rect 2065 2746 2071 2748
rect 2127 2746 2151 2748
rect 2207 2746 2231 2748
rect 2287 2746 2311 2748
rect 2367 2746 2373 2748
rect 2127 2694 2129 2746
rect 2309 2694 2311 2746
rect 2065 2692 2071 2694
rect 2127 2692 2151 2694
rect 2207 2692 2231 2694
rect 2287 2692 2311 2694
rect 2367 2692 2373 2694
rect 2065 2683 2373 2692
rect 2516 2446 2544 3878
rect 3528 3398 3556 3878
rect 3804 3670 3832 4082
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3896 3602 3924 4558
rect 3988 4146 4016 5766
rect 4172 5681 4200 6666
rect 4264 6254 4292 6938
rect 4632 6934 4660 7414
rect 4724 7398 4936 7426
rect 5356 7414 5408 7420
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4356 6458 4384 6734
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4356 6118 4384 6258
rect 4448 6186 4476 6734
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 6458 4568 6598
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4526 6352 4582 6361
rect 4526 6287 4528 6296
rect 4580 6287 4582 6296
rect 4528 6258 4580 6264
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4296 6012 4604 6021
rect 4296 6010 4302 6012
rect 4358 6010 4382 6012
rect 4438 6010 4462 6012
rect 4518 6010 4542 6012
rect 4598 6010 4604 6012
rect 4358 5958 4360 6010
rect 4540 5958 4542 6010
rect 4296 5956 4302 5958
rect 4358 5956 4382 5958
rect 4438 5956 4462 5958
rect 4518 5956 4542 5958
rect 4598 5956 4604 5958
rect 4296 5947 4604 5956
rect 4158 5672 4214 5681
rect 4158 5607 4214 5616
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4172 4162 4200 5510
rect 4264 5370 4292 5510
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4296 4924 4604 4933
rect 4296 4922 4302 4924
rect 4358 4922 4382 4924
rect 4438 4922 4462 4924
rect 4518 4922 4542 4924
rect 4598 4922 4604 4924
rect 4358 4870 4360 4922
rect 4540 4870 4542 4922
rect 4296 4868 4302 4870
rect 4358 4868 4382 4870
rect 4438 4868 4462 4870
rect 4518 4868 4542 4870
rect 4598 4868 4604 4870
rect 4296 4859 4604 4868
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4282 4476 4490
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4080 4134 4200 4162
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 2725 3292 3033 3301
rect 2725 3290 2731 3292
rect 2787 3290 2811 3292
rect 2867 3290 2891 3292
rect 2947 3290 2971 3292
rect 3027 3290 3033 3292
rect 2787 3238 2789 3290
rect 2969 3238 2971 3290
rect 2725 3236 2731 3238
rect 2787 3236 2811 3238
rect 2867 3236 2891 3238
rect 2947 3236 2971 3238
rect 3027 3236 3033 3238
rect 2725 3227 3033 3236
rect 3896 3194 3924 3538
rect 3988 3516 4016 4082
rect 4080 3618 4108 4134
rect 4540 4078 4568 4558
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4172 3738 4200 4014
rect 4296 3836 4604 3845
rect 4296 3834 4302 3836
rect 4358 3834 4382 3836
rect 4438 3834 4462 3836
rect 4518 3834 4542 3836
rect 4598 3834 4604 3836
rect 4358 3782 4360 3834
rect 4540 3782 4542 3834
rect 4296 3780 4302 3782
rect 4358 3780 4382 3782
rect 4438 3780 4462 3782
rect 4518 3780 4542 3782
rect 4598 3780 4604 3782
rect 4296 3771 4604 3780
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4080 3590 4292 3618
rect 4068 3528 4120 3534
rect 3988 3488 4068 3516
rect 4068 3470 4120 3476
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 4080 2514 4108 3470
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 4172 2650 4200 3402
rect 4264 2854 4292 3590
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4448 3058 4476 3334
rect 4540 3194 4568 3334
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4632 3126 4660 6870
rect 4724 6458 4752 7278
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4724 6118 4752 6258
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4724 3534 4752 5510
rect 4816 4622 4844 7142
rect 4908 7002 4936 7398
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 5000 6798 5028 7142
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4956 6556 5264 6565
rect 4956 6554 4962 6556
rect 5018 6554 5042 6556
rect 5098 6554 5122 6556
rect 5178 6554 5202 6556
rect 5258 6554 5264 6556
rect 5018 6502 5020 6554
rect 5200 6502 5202 6554
rect 4956 6500 4962 6502
rect 5018 6500 5042 6502
rect 5098 6500 5122 6502
rect 5178 6500 5202 6502
rect 5258 6500 5264 6502
rect 4956 6491 5264 6500
rect 5368 6322 5396 7414
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6662 5488 7346
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4908 5914 4936 6190
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5000 5642 5028 6054
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 5092 5556 5120 6258
rect 5460 6254 5488 6598
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5172 5568 5224 5574
rect 5092 5528 5172 5556
rect 5172 5510 5224 5516
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 4956 5468 5264 5477
rect 4956 5466 4962 5468
rect 5018 5466 5042 5468
rect 5098 5466 5122 5468
rect 5178 5466 5202 5468
rect 5258 5466 5264 5468
rect 5018 5414 5020 5466
rect 5200 5414 5202 5466
rect 4956 5412 4962 5414
rect 5018 5412 5042 5414
rect 5098 5412 5122 5414
rect 5178 5412 5202 5414
rect 5258 5412 5264 5414
rect 4956 5403 5264 5412
rect 5368 5234 5396 5510
rect 5460 5386 5488 6190
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5460 5358 5580 5386
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5092 4826 5120 4966
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5092 4622 5120 4762
rect 5184 4690 5212 4966
rect 5276 4690 5304 5034
rect 5368 5012 5396 5170
rect 5448 5024 5500 5030
rect 5368 4984 5448 5012
rect 5552 5012 5580 5358
rect 5644 5166 5672 5510
rect 5736 5234 5764 6054
rect 5920 5710 5948 7822
rect 6104 7750 6132 8026
rect 6368 7880 6420 7886
rect 6196 7840 6368 7868
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5552 4984 5672 5012
rect 5448 4966 5500 4972
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5184 4570 5212 4626
rect 5460 4570 5488 4626
rect 5184 4542 5396 4570
rect 5460 4542 5580 4570
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 3534 4844 4422
rect 4956 4380 5264 4389
rect 4956 4378 4962 4380
rect 5018 4378 5042 4380
rect 5098 4378 5122 4380
rect 5178 4378 5202 4380
rect 5258 4378 5264 4380
rect 5018 4326 5020 4378
rect 5200 4326 5202 4378
rect 4956 4324 4962 4326
rect 5018 4324 5042 4326
rect 5098 4324 5122 4326
rect 5178 4324 5202 4326
rect 5258 4324 5264 4326
rect 4956 4315 5264 4324
rect 5368 4282 5396 4542
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4162 5488 4422
rect 5552 4282 5580 4542
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5368 4146 5488 4162
rect 5356 4140 5488 4146
rect 5408 4134 5488 4140
rect 5356 4082 5408 4088
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 4908 3738 4936 3878
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4908 3466 4936 3674
rect 5092 3534 5120 3878
rect 5276 3534 5304 3878
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5552 3534 5580 3606
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4956 3292 5264 3301
rect 4956 3290 4962 3292
rect 5018 3290 5042 3292
rect 5098 3290 5122 3292
rect 5178 3290 5202 3292
rect 5258 3290 5264 3292
rect 5018 3238 5020 3290
rect 5200 3238 5202 3290
rect 4956 3236 4962 3238
rect 5018 3236 5042 3238
rect 5098 3236 5122 3238
rect 5178 3236 5202 3238
rect 5258 3236 5264 3238
rect 4956 3227 5264 3236
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4296 2748 4604 2757
rect 4296 2746 4302 2748
rect 4358 2746 4382 2748
rect 4438 2746 4462 2748
rect 4518 2746 4542 2748
rect 4598 2746 4604 2748
rect 4358 2694 4360 2746
rect 4540 2694 4542 2746
rect 4296 2692 4302 2694
rect 4358 2692 4382 2694
rect 4438 2692 4462 2694
rect 4518 2692 4542 2694
rect 4598 2692 4604 2694
rect 4296 2683 4604 2692
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4724 2446 4752 2790
rect 5552 2650 5580 2994
rect 5644 2854 5672 4984
rect 5920 4826 5948 5646
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5920 4282 5948 4762
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 6012 4146 6040 4694
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5736 3126 5764 3470
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 6012 3058 6040 4082
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 2446 5672 2790
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2504 2440 2556 2446
rect 4712 2440 4764 2446
rect 2504 2382 2556 2388
rect 2608 2378 2820 2394
rect 4712 2382 4764 2388
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 2608 2372 2832 2378
rect 2608 2366 2780 2372
rect 1490 1592 1546 1601
rect 1490 1527 1546 1536
rect 2608 800 2636 2366
rect 2780 2314 2832 2320
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 2725 2204 3033 2213
rect 2725 2202 2731 2204
rect 2787 2202 2811 2204
rect 2867 2202 2891 2204
rect 2947 2202 2971 2204
rect 3027 2202 3033 2204
rect 2787 2150 2789 2202
rect 2969 2150 2971 2202
rect 2725 2148 2731 2150
rect 2787 2148 2811 2150
rect 2867 2148 2891 2150
rect 2947 2148 2971 2150
rect 3027 2148 3033 2150
rect 2725 2139 3033 2148
rect 4540 800 4568 2314
rect 6196 2310 6224 7840
rect 6368 7822 6420 7828
rect 6828 7880 6880 7886
rect 6932 7868 6960 9318
rect 7012 7948 7064 7954
rect 7116 7936 7144 9318
rect 7187 8732 7495 8741
rect 7187 8730 7193 8732
rect 7249 8730 7273 8732
rect 7329 8730 7353 8732
rect 7409 8730 7433 8732
rect 7489 8730 7495 8732
rect 7249 8678 7251 8730
rect 7431 8678 7433 8730
rect 7187 8676 7193 8678
rect 7249 8676 7273 8678
rect 7329 8676 7353 8678
rect 7409 8676 7433 8678
rect 7489 8676 7495 8678
rect 7187 8667 7495 8676
rect 7196 7948 7248 7954
rect 7116 7908 7196 7936
rect 7012 7890 7064 7896
rect 7196 7890 7248 7896
rect 6880 7840 6960 7868
rect 6828 7822 6880 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 6798 6316 7686
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6380 6458 6408 7346
rect 6840 7274 6868 7822
rect 7024 7750 7052 7890
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7546 7052 7686
rect 7187 7644 7495 7653
rect 7187 7642 7193 7644
rect 7249 7642 7273 7644
rect 7329 7642 7353 7644
rect 7409 7642 7433 7644
rect 7489 7642 7495 7644
rect 7249 7590 7251 7642
rect 7431 7590 7433 7642
rect 7187 7588 7193 7590
rect 7249 7588 7273 7590
rect 7329 7588 7353 7590
rect 7409 7588 7433 7590
rect 7489 7588 7495 7590
rect 7187 7579 7495 7588
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6527 7100 6835 7109
rect 6527 7098 6533 7100
rect 6589 7098 6613 7100
rect 6669 7098 6693 7100
rect 6749 7098 6773 7100
rect 6829 7098 6835 7100
rect 6589 7046 6591 7098
rect 6771 7046 6773 7098
rect 6527 7044 6533 7046
rect 6589 7044 6613 7046
rect 6669 7044 6693 7046
rect 6749 7044 6773 7046
rect 6829 7044 6835 7046
rect 6527 7035 6835 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6527 6012 6835 6021
rect 6527 6010 6533 6012
rect 6589 6010 6613 6012
rect 6669 6010 6693 6012
rect 6749 6010 6773 6012
rect 6829 6010 6835 6012
rect 6589 5958 6591 6010
rect 6771 5958 6773 6010
rect 6527 5956 6533 5958
rect 6589 5956 6613 5958
rect 6669 5956 6693 5958
rect 6749 5956 6773 5958
rect 6829 5956 6835 5958
rect 6527 5947 6835 5956
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6288 5370 6316 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6564 5030 6592 5646
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5302 6868 5510
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 4282 6316 4490
rect 6380 4282 6408 4966
rect 6527 4924 6835 4933
rect 6527 4922 6533 4924
rect 6589 4922 6613 4924
rect 6669 4922 6693 4924
rect 6749 4922 6773 4924
rect 6829 4922 6835 4924
rect 6589 4870 6591 4922
rect 6771 4870 6773 4922
rect 6527 4868 6533 4870
rect 6589 4868 6613 4870
rect 6669 4868 6693 4870
rect 6749 4868 6773 4870
rect 6829 4868 6835 4870
rect 6527 4859 6835 4868
rect 6932 4434 6960 6802
rect 7024 6458 7052 7482
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7116 7002 7144 7142
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7208 6644 7236 7142
rect 7484 6798 7512 7414
rect 7668 7410 7696 9454
rect 7944 9178 7972 9930
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7852 8634 7880 9114
rect 8036 8974 8064 9862
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8128 9178 8156 9522
rect 8220 9382 8248 10639
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 9048 10554 9076 12534
rect 9402 12336 9458 12345
rect 9324 12294 9402 12322
rect 9324 10810 9352 12294
rect 9402 12271 9458 12280
rect 9418 10908 9726 10917
rect 9418 10906 9424 10908
rect 9480 10906 9504 10908
rect 9560 10906 9584 10908
rect 9640 10906 9664 10908
rect 9720 10906 9726 10908
rect 9480 10854 9482 10906
rect 9662 10854 9664 10906
rect 9418 10852 9424 10854
rect 9480 10852 9504 10854
rect 9560 10852 9584 10854
rect 9640 10852 9664 10854
rect 9720 10852 9726 10854
rect 9418 10843 9726 10852
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 8404 9926 8432 10542
rect 9048 10526 9260 10554
rect 8758 10364 9066 10373
rect 8758 10362 8764 10364
rect 8820 10362 8844 10364
rect 8900 10362 8924 10364
rect 8980 10362 9004 10364
rect 9060 10362 9066 10364
rect 8820 10310 8822 10362
rect 9002 10310 9004 10362
rect 8758 10308 8764 10310
rect 8820 10308 8844 10310
rect 8900 10308 8924 10310
rect 8980 10308 9004 10310
rect 9060 10308 9066 10310
rect 8758 10299 9066 10308
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8404 9654 8432 9862
rect 8956 9654 8984 9862
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8312 9042 8340 9454
rect 8758 9276 9066 9285
rect 8758 9274 8764 9276
rect 8820 9274 8844 9276
rect 8900 9274 8924 9276
rect 8980 9274 9004 9276
rect 9060 9274 9066 9276
rect 8820 9222 8822 9274
rect 9002 9222 9004 9274
rect 8758 9220 8764 9222
rect 8820 9220 8844 9222
rect 8900 9220 8924 9222
rect 8980 9220 9004 9222
rect 9060 9220 9066 9222
rect 8758 9211 9066 9220
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7576 6730 7604 7278
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7116 6616 7236 6644
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 5574 7052 6122
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7116 5370 7144 6616
rect 7187 6556 7495 6565
rect 7187 6554 7193 6556
rect 7249 6554 7273 6556
rect 7329 6554 7353 6556
rect 7409 6554 7433 6556
rect 7489 6554 7495 6556
rect 7249 6502 7251 6554
rect 7431 6502 7433 6554
rect 7187 6500 7193 6502
rect 7249 6500 7273 6502
rect 7329 6500 7353 6502
rect 7409 6500 7433 6502
rect 7489 6500 7495 6502
rect 7187 6491 7495 6500
rect 7576 6458 7604 6666
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7668 6338 7696 7210
rect 7760 7002 7788 7958
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7576 6310 7696 6338
rect 7576 5710 7604 6310
rect 7852 6254 7880 8570
rect 7944 8294 7972 8842
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7546 7972 8230
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 7002 8064 7346
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7187 5468 7495 5477
rect 7187 5466 7193 5468
rect 7249 5466 7273 5468
rect 7329 5466 7353 5468
rect 7409 5466 7433 5468
rect 7489 5466 7495 5468
rect 7249 5414 7251 5466
rect 7431 5414 7433 5466
rect 7187 5412 7193 5414
rect 7249 5412 7273 5414
rect 7329 5412 7353 5414
rect 7409 5412 7433 5414
rect 7489 5412 7495 5414
rect 7187 5403 7495 5412
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 7024 4554 7052 5306
rect 7116 4554 7144 5306
rect 7852 5234 7880 5850
rect 7944 5234 7972 6190
rect 8036 5914 8064 6802
rect 8128 6458 8156 7822
rect 8312 7410 8340 8978
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8220 6390 8248 7142
rect 8404 7002 8432 7346
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5302 8064 5510
rect 8496 5302 8524 8774
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7300 4622 7328 5102
rect 7392 4690 7420 5102
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6932 4406 7144 4434
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6288 4078 6316 4218
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6288 3534 6316 4014
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6288 3058 6316 3470
rect 6380 3058 6408 3946
rect 6527 3836 6835 3845
rect 6527 3834 6533 3836
rect 6589 3834 6613 3836
rect 6669 3834 6693 3836
rect 6749 3834 6773 3836
rect 6829 3834 6835 3836
rect 6589 3782 6591 3834
rect 6771 3782 6773 3834
rect 6527 3780 6533 3782
rect 6589 3780 6613 3782
rect 6669 3780 6693 3782
rect 6749 3780 6773 3782
rect 6829 3780 6835 3782
rect 6527 3771 6835 3780
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 3194 6960 3470
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7024 3058 7052 4218
rect 7116 4146 7144 4406
rect 7187 4380 7495 4389
rect 7187 4378 7193 4380
rect 7249 4378 7273 4380
rect 7329 4378 7353 4380
rect 7409 4378 7433 4380
rect 7489 4378 7495 4380
rect 7249 4326 7251 4378
rect 7431 4326 7433 4378
rect 7187 4324 7193 4326
rect 7249 4324 7273 4326
rect 7329 4324 7353 4326
rect 7409 4324 7433 4326
rect 7489 4324 7495 4326
rect 7187 4315 7495 4324
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7116 3058 7144 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3738 7328 3878
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7187 3292 7495 3301
rect 7187 3290 7193 3292
rect 7249 3290 7273 3292
rect 7329 3290 7353 3292
rect 7409 3290 7433 3292
rect 7489 3290 7495 3292
rect 7249 3238 7251 3290
rect 7431 3238 7433 3290
rect 7187 3236 7193 3238
rect 7249 3236 7273 3238
rect 7329 3236 7353 3238
rect 7409 3236 7433 3238
rect 7489 3236 7495 3238
rect 7187 3227 7495 3236
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7208 3058 7236 3130
rect 7576 3058 7604 3334
rect 7852 3194 7880 5170
rect 7944 4146 7972 5170
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4282 8340 4966
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 3058 7972 4082
rect 8588 3466 8616 8978
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8430 9168 9998
rect 9232 8634 9260 10526
rect 10336 10266 10364 12534
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9418 9820 9726 9829
rect 9418 9818 9424 9820
rect 9480 9818 9504 9820
rect 9560 9818 9584 9820
rect 9640 9818 9664 9820
rect 9720 9818 9726 9820
rect 9480 9766 9482 9818
rect 9662 9766 9664 9818
rect 9418 9764 9424 9766
rect 9480 9764 9504 9766
rect 9560 9764 9584 9766
rect 9640 9764 9664 9766
rect 9720 9764 9726 9766
rect 9418 9755 9726 9764
rect 9784 9450 9812 9930
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9784 9042 9812 9386
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9678 8936 9734 8945
rect 9678 8871 9680 8880
rect 9732 8871 9734 8880
rect 9680 8842 9732 8848
rect 9418 8732 9726 8741
rect 9418 8730 9424 8732
rect 9480 8730 9504 8732
rect 9560 8730 9584 8732
rect 9640 8730 9664 8732
rect 9720 8730 9726 8732
rect 9480 8678 9482 8730
rect 9662 8678 9664 8730
rect 9418 8676 9424 8678
rect 9480 8676 9504 8678
rect 9560 8676 9584 8678
rect 9640 8676 9664 8678
rect 9720 8676 9726 8678
rect 9418 8667 9726 8676
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8758 8188 9066 8197
rect 8758 8186 8764 8188
rect 8820 8186 8844 8188
rect 8900 8186 8924 8188
rect 8980 8186 9004 8188
rect 9060 8186 9066 8188
rect 8820 8134 8822 8186
rect 9002 8134 9004 8186
rect 8758 8132 8764 8134
rect 8820 8132 8844 8134
rect 8900 8132 8924 8134
rect 8980 8132 9004 8134
rect 9060 8132 9066 8134
rect 8758 8123 9066 8132
rect 8758 7100 9066 7109
rect 8758 7098 8764 7100
rect 8820 7098 8844 7100
rect 8900 7098 8924 7100
rect 8980 7098 9004 7100
rect 9060 7098 9066 7100
rect 8820 7046 8822 7098
rect 9002 7046 9004 7098
rect 8758 7044 8764 7046
rect 8820 7044 8844 7046
rect 8900 7044 8924 7046
rect 8980 7044 9004 7046
rect 9060 7044 9066 7046
rect 8758 7035 9066 7044
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8772 6458 8800 6802
rect 9324 6458 9352 8434
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9418 7644 9726 7653
rect 9418 7642 9424 7644
rect 9480 7642 9504 7644
rect 9560 7642 9584 7644
rect 9640 7642 9664 7644
rect 9720 7642 9726 7644
rect 9480 7590 9482 7642
rect 9662 7590 9664 7642
rect 9418 7588 9424 7590
rect 9480 7588 9504 7590
rect 9560 7588 9584 7590
rect 9640 7588 9664 7590
rect 9720 7588 9726 7590
rect 9418 7579 9726 7588
rect 9968 7585 9996 7686
rect 9954 7576 10010 7585
rect 9954 7511 10010 7520
rect 9418 6556 9726 6565
rect 9418 6554 9424 6556
rect 9480 6554 9504 6556
rect 9560 6554 9584 6556
rect 9640 6554 9664 6556
rect 9720 6554 9726 6556
rect 9480 6502 9482 6554
rect 9662 6502 9664 6554
rect 9418 6500 9424 6502
rect 9480 6500 9504 6502
rect 9560 6500 9584 6502
rect 9640 6500 9664 6502
rect 9720 6500 9726 6502
rect 9418 6491 9726 6500
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8758 6012 9066 6021
rect 8758 6010 8764 6012
rect 8820 6010 8844 6012
rect 8900 6010 8924 6012
rect 8980 6010 9004 6012
rect 9060 6010 9066 6012
rect 8820 5958 8822 6010
rect 9002 5958 9004 6010
rect 8758 5956 8764 5958
rect 8820 5956 8844 5958
rect 8900 5956 8924 5958
rect 8980 5956 9004 5958
rect 9060 5956 9066 5958
rect 8758 5947 9066 5956
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9324 5370 9352 5782
rect 10046 5536 10102 5545
rect 9418 5468 9726 5477
rect 10046 5471 10102 5480
rect 9418 5466 9424 5468
rect 9480 5466 9504 5468
rect 9560 5466 9584 5468
rect 9640 5466 9664 5468
rect 9720 5466 9726 5468
rect 9480 5414 9482 5466
rect 9662 5414 9664 5466
rect 9418 5412 9424 5414
rect 9480 5412 9504 5414
rect 9560 5412 9584 5414
rect 9640 5412 9664 5414
rect 9720 5412 9726 5414
rect 9418 5403 9726 5412
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 8758 4924 9066 4933
rect 8758 4922 8764 4924
rect 8820 4922 8844 4924
rect 8900 4922 8924 4924
rect 8980 4922 9004 4924
rect 9060 4922 9066 4924
rect 8820 4870 8822 4922
rect 9002 4870 9004 4922
rect 8758 4868 8764 4870
rect 8820 4868 8844 4870
rect 8900 4868 8924 4870
rect 8980 4868 9004 4870
rect 9060 4868 9066 4870
rect 8758 4859 9066 4868
rect 8758 3836 9066 3845
rect 8758 3834 8764 3836
rect 8820 3834 8844 3836
rect 8900 3834 8924 3836
rect 8980 3834 9004 3836
rect 9060 3834 9066 3836
rect 8820 3782 8822 3834
rect 9002 3782 9004 3834
rect 8758 3780 8764 3782
rect 8820 3780 8844 3782
rect 8900 3780 8924 3782
rect 8980 3780 9004 3782
rect 9060 3780 9066 3782
rect 8758 3771 9066 3780
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 6527 2748 6835 2757
rect 6527 2746 6533 2748
rect 6589 2746 6613 2748
rect 6669 2746 6693 2748
rect 6749 2746 6773 2748
rect 6829 2746 6835 2748
rect 6589 2694 6591 2746
rect 6771 2694 6773 2746
rect 6527 2692 6533 2694
rect 6589 2692 6613 2694
rect 6669 2692 6693 2694
rect 6749 2692 6773 2694
rect 6829 2692 6835 2694
rect 6527 2683 6835 2692
rect 7208 2446 7236 2790
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 8220 2378 8248 2790
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 4956 2204 5264 2213
rect 4956 2202 4962 2204
rect 5018 2202 5042 2204
rect 5098 2202 5122 2204
rect 5178 2202 5202 2204
rect 5258 2202 5264 2204
rect 5018 2150 5020 2202
rect 5200 2150 5202 2202
rect 4956 2148 4962 2150
rect 5018 2148 5042 2150
rect 5098 2148 5122 2150
rect 5178 2148 5202 2150
rect 5258 2148 5264 2150
rect 4956 2139 5264 2148
rect 5828 800 5856 2246
rect 7187 2204 7495 2213
rect 7187 2202 7193 2204
rect 7249 2202 7273 2204
rect 7329 2202 7353 2204
rect 7409 2202 7433 2204
rect 7489 2202 7495 2204
rect 7249 2150 7251 2202
rect 7431 2150 7433 2202
rect 7187 2148 7193 2150
rect 7249 2148 7273 2150
rect 7329 2148 7353 2150
rect 7409 2148 7433 2150
rect 7489 2148 7495 2150
rect 7187 2139 7495 2148
rect 7760 800 7788 2246
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 8680 785 8708 3334
rect 9048 2854 9076 3470
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8758 2748 9066 2757
rect 8758 2746 8764 2748
rect 8820 2746 8844 2748
rect 8900 2746 8924 2748
rect 8980 2746 9004 2748
rect 9060 2746 9066 2748
rect 8820 2694 8822 2746
rect 9002 2694 9004 2746
rect 8758 2692 8764 2694
rect 8820 2692 8844 2694
rect 8900 2692 8924 2694
rect 8980 2692 9004 2694
rect 9060 2692 9066 2694
rect 8758 2683 9066 2692
rect 9324 2446 9352 5306
rect 10060 5302 10088 5471
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9418 4380 9726 4389
rect 9418 4378 9424 4380
rect 9480 4378 9504 4380
rect 9560 4378 9584 4380
rect 9640 4378 9664 4380
rect 9720 4378 9726 4380
rect 9480 4326 9482 4378
rect 9662 4326 9664 4378
rect 9418 4324 9424 4326
rect 9480 4324 9504 4326
rect 9560 4324 9584 4326
rect 9640 4324 9664 4326
rect 9720 4324 9726 4326
rect 9418 4315 9726 4324
rect 9784 4282 9812 4558
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9876 4185 9904 4422
rect 9862 4176 9918 4185
rect 9862 4111 9918 4120
rect 9418 3292 9726 3301
rect 9418 3290 9424 3292
rect 9480 3290 9504 3292
rect 9560 3290 9584 3292
rect 9640 3290 9664 3292
rect 9720 3290 9726 3292
rect 9480 3238 9482 3290
rect 9662 3238 9664 3290
rect 9418 3236 9424 3238
rect 9480 3236 9504 3238
rect 9560 3236 9584 3238
rect 9640 3236 9664 3238
rect 9720 3236 9726 3238
rect 9418 3227 9726 3236
rect 9772 2848 9824 2854
rect 9770 2816 9772 2825
rect 9824 2816 9826 2825
rect 9770 2751 9826 2760
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 800 9076 2246
rect 9418 2204 9726 2213
rect 9418 2202 9424 2204
rect 9480 2202 9504 2204
rect 9560 2202 9584 2204
rect 9640 2202 9664 2204
rect 9720 2202 9726 2204
rect 9480 2150 9482 2202
rect 9662 2150 9664 2202
rect 9418 2148 9424 2150
rect 9480 2148 9504 2150
rect 9560 2148 9584 2150
rect 9640 2148 9664 2150
rect 9720 2148 9726 2150
rect 9418 2139 9726 2148
rect 10980 800 11008 2450
rect 8666 776 8722 785
rect 8666 711 8722 720
rect 9034 0 9090 800
rect 10966 0 11022 800
<< via2 >>
rect 3054 12960 3110 13016
rect 1582 11600 1638 11656
rect 2731 10906 2787 10908
rect 2811 10906 2867 10908
rect 2891 10906 2947 10908
rect 2971 10906 3027 10908
rect 2731 10854 2777 10906
rect 2777 10854 2787 10906
rect 2811 10854 2841 10906
rect 2841 10854 2853 10906
rect 2853 10854 2867 10906
rect 2891 10854 2905 10906
rect 2905 10854 2917 10906
rect 2917 10854 2947 10906
rect 2971 10854 2981 10906
rect 2981 10854 3027 10906
rect 2731 10852 2787 10854
rect 2811 10852 2867 10854
rect 2891 10852 2947 10854
rect 2971 10852 3027 10854
rect 4962 10906 5018 10908
rect 5042 10906 5098 10908
rect 5122 10906 5178 10908
rect 5202 10906 5258 10908
rect 4962 10854 5008 10906
rect 5008 10854 5018 10906
rect 5042 10854 5072 10906
rect 5072 10854 5084 10906
rect 5084 10854 5098 10906
rect 5122 10854 5136 10906
rect 5136 10854 5148 10906
rect 5148 10854 5178 10906
rect 5202 10854 5212 10906
rect 5212 10854 5258 10906
rect 4962 10852 5018 10854
rect 5042 10852 5098 10854
rect 5122 10852 5178 10854
rect 5202 10852 5258 10854
rect 7193 10906 7249 10908
rect 7273 10906 7329 10908
rect 7353 10906 7409 10908
rect 7433 10906 7489 10908
rect 7193 10854 7239 10906
rect 7239 10854 7249 10906
rect 7273 10854 7303 10906
rect 7303 10854 7315 10906
rect 7315 10854 7329 10906
rect 7353 10854 7367 10906
rect 7367 10854 7379 10906
rect 7379 10854 7409 10906
rect 7433 10854 7443 10906
rect 7443 10854 7489 10906
rect 7193 10852 7249 10854
rect 7273 10852 7329 10854
rect 7353 10852 7409 10854
rect 7433 10852 7489 10854
rect 8206 10648 8262 10704
rect 2071 10362 2127 10364
rect 2151 10362 2207 10364
rect 2231 10362 2287 10364
rect 2311 10362 2367 10364
rect 2071 10310 2117 10362
rect 2117 10310 2127 10362
rect 2151 10310 2181 10362
rect 2181 10310 2193 10362
rect 2193 10310 2207 10362
rect 2231 10310 2245 10362
rect 2245 10310 2257 10362
rect 2257 10310 2287 10362
rect 2311 10310 2321 10362
rect 2321 10310 2367 10362
rect 2071 10308 2127 10310
rect 2151 10308 2207 10310
rect 2231 10308 2287 10310
rect 2311 10308 2367 10310
rect 1490 9560 1546 9616
rect 2071 9274 2127 9276
rect 2151 9274 2207 9276
rect 2231 9274 2287 9276
rect 2311 9274 2367 9276
rect 2071 9222 2117 9274
rect 2117 9222 2127 9274
rect 2151 9222 2181 9274
rect 2181 9222 2193 9274
rect 2193 9222 2207 9274
rect 2231 9222 2245 9274
rect 2245 9222 2257 9274
rect 2257 9222 2287 9274
rect 2311 9222 2321 9274
rect 2321 9222 2367 9274
rect 2071 9220 2127 9222
rect 2151 9220 2207 9222
rect 2231 9220 2287 9222
rect 2311 9220 2367 9222
rect 938 8200 994 8256
rect 2071 8186 2127 8188
rect 2151 8186 2207 8188
rect 2231 8186 2287 8188
rect 2311 8186 2367 8188
rect 2071 8134 2117 8186
rect 2117 8134 2127 8186
rect 2151 8134 2181 8186
rect 2181 8134 2193 8186
rect 2193 8134 2207 8186
rect 2231 8134 2245 8186
rect 2245 8134 2257 8186
rect 2257 8134 2287 8186
rect 2311 8134 2321 8186
rect 2321 8134 2367 8186
rect 2071 8132 2127 8134
rect 2151 8132 2207 8134
rect 2231 8132 2287 8134
rect 2311 8132 2367 8134
rect 2071 7098 2127 7100
rect 2151 7098 2207 7100
rect 2231 7098 2287 7100
rect 2311 7098 2367 7100
rect 2071 7046 2117 7098
rect 2117 7046 2127 7098
rect 2151 7046 2181 7098
rect 2181 7046 2193 7098
rect 2193 7046 2207 7098
rect 2231 7046 2245 7098
rect 2245 7046 2257 7098
rect 2257 7046 2287 7098
rect 2311 7046 2321 7098
rect 2321 7046 2367 7098
rect 2071 7044 2127 7046
rect 2151 7044 2207 7046
rect 2231 7044 2287 7046
rect 2311 7044 2367 7046
rect 2731 9818 2787 9820
rect 2811 9818 2867 9820
rect 2891 9818 2947 9820
rect 2971 9818 3027 9820
rect 2731 9766 2777 9818
rect 2777 9766 2787 9818
rect 2811 9766 2841 9818
rect 2841 9766 2853 9818
rect 2853 9766 2867 9818
rect 2891 9766 2905 9818
rect 2905 9766 2917 9818
rect 2917 9766 2947 9818
rect 2971 9766 2981 9818
rect 2981 9766 3027 9818
rect 2731 9764 2787 9766
rect 2811 9764 2867 9766
rect 2891 9764 2947 9766
rect 2971 9764 3027 9766
rect 4302 10362 4358 10364
rect 4382 10362 4438 10364
rect 4462 10362 4518 10364
rect 4542 10362 4598 10364
rect 4302 10310 4348 10362
rect 4348 10310 4358 10362
rect 4382 10310 4412 10362
rect 4412 10310 4424 10362
rect 4424 10310 4438 10362
rect 4462 10310 4476 10362
rect 4476 10310 4488 10362
rect 4488 10310 4518 10362
rect 4542 10310 4552 10362
rect 4552 10310 4598 10362
rect 4302 10308 4358 10310
rect 4382 10308 4438 10310
rect 4462 10308 4518 10310
rect 4542 10308 4598 10310
rect 2731 8730 2787 8732
rect 2811 8730 2867 8732
rect 2891 8730 2947 8732
rect 2971 8730 3027 8732
rect 2731 8678 2777 8730
rect 2777 8678 2787 8730
rect 2811 8678 2841 8730
rect 2841 8678 2853 8730
rect 2853 8678 2867 8730
rect 2891 8678 2905 8730
rect 2905 8678 2917 8730
rect 2917 8678 2947 8730
rect 2971 8678 2981 8730
rect 2981 8678 3027 8730
rect 2731 8676 2787 8678
rect 2811 8676 2867 8678
rect 2891 8676 2947 8678
rect 2971 8676 3027 8678
rect 2731 7642 2787 7644
rect 2811 7642 2867 7644
rect 2891 7642 2947 7644
rect 2971 7642 3027 7644
rect 2731 7590 2777 7642
rect 2777 7590 2787 7642
rect 2811 7590 2841 7642
rect 2841 7590 2853 7642
rect 2853 7590 2867 7642
rect 2891 7590 2905 7642
rect 2905 7590 2917 7642
rect 2917 7590 2947 7642
rect 2971 7590 2981 7642
rect 2981 7590 3027 7642
rect 2731 7588 2787 7590
rect 2811 7588 2867 7590
rect 2891 7588 2947 7590
rect 2971 7588 3027 7590
rect 4302 9274 4358 9276
rect 4382 9274 4438 9276
rect 4462 9274 4518 9276
rect 4542 9274 4598 9276
rect 4302 9222 4348 9274
rect 4348 9222 4358 9274
rect 4382 9222 4412 9274
rect 4412 9222 4424 9274
rect 4424 9222 4438 9274
rect 4462 9222 4476 9274
rect 4476 9222 4488 9274
rect 4488 9222 4518 9274
rect 4542 9222 4552 9274
rect 4552 9222 4598 9274
rect 4302 9220 4358 9222
rect 4382 9220 4438 9222
rect 4462 9220 4518 9222
rect 4542 9220 4598 9222
rect 6533 10362 6589 10364
rect 6613 10362 6669 10364
rect 6693 10362 6749 10364
rect 6773 10362 6829 10364
rect 6533 10310 6579 10362
rect 6579 10310 6589 10362
rect 6613 10310 6643 10362
rect 6643 10310 6655 10362
rect 6655 10310 6669 10362
rect 6693 10310 6707 10362
rect 6707 10310 6719 10362
rect 6719 10310 6749 10362
rect 6773 10310 6783 10362
rect 6783 10310 6829 10362
rect 6533 10308 6589 10310
rect 6613 10308 6669 10310
rect 6693 10308 6749 10310
rect 6773 10308 6829 10310
rect 4962 9818 5018 9820
rect 5042 9818 5098 9820
rect 5122 9818 5178 9820
rect 5202 9818 5258 9820
rect 4962 9766 5008 9818
rect 5008 9766 5018 9818
rect 5042 9766 5072 9818
rect 5072 9766 5084 9818
rect 5084 9766 5098 9818
rect 5122 9766 5136 9818
rect 5136 9766 5148 9818
rect 5148 9766 5178 9818
rect 5202 9766 5212 9818
rect 5212 9766 5258 9818
rect 4962 9764 5018 9766
rect 5042 9764 5098 9766
rect 5122 9764 5178 9766
rect 5202 9764 5258 9766
rect 4962 8730 5018 8732
rect 5042 8730 5098 8732
rect 5122 8730 5178 8732
rect 5202 8730 5258 8732
rect 4962 8678 5008 8730
rect 5008 8678 5018 8730
rect 5042 8678 5072 8730
rect 5072 8678 5084 8730
rect 5084 8678 5098 8730
rect 5122 8678 5136 8730
rect 5136 8678 5148 8730
rect 5148 8678 5178 8730
rect 5202 8678 5212 8730
rect 5212 8678 5258 8730
rect 4962 8676 5018 8678
rect 5042 8676 5098 8678
rect 5122 8676 5178 8678
rect 5202 8676 5258 8678
rect 7193 9818 7249 9820
rect 7273 9818 7329 9820
rect 7353 9818 7409 9820
rect 7433 9818 7489 9820
rect 7193 9766 7239 9818
rect 7239 9766 7249 9818
rect 7273 9766 7303 9818
rect 7303 9766 7315 9818
rect 7315 9766 7329 9818
rect 7353 9766 7367 9818
rect 7367 9766 7379 9818
rect 7379 9766 7409 9818
rect 7433 9766 7443 9818
rect 7443 9766 7489 9818
rect 7193 9764 7249 9766
rect 7273 9764 7329 9766
rect 7353 9764 7409 9766
rect 7433 9764 7489 9766
rect 6533 9274 6589 9276
rect 6613 9274 6669 9276
rect 6693 9274 6749 9276
rect 6773 9274 6829 9276
rect 6533 9222 6579 9274
rect 6579 9222 6589 9274
rect 6613 9222 6643 9274
rect 6643 9222 6655 9274
rect 6655 9222 6669 9274
rect 6693 9222 6707 9274
rect 6707 9222 6719 9274
rect 6719 9222 6749 9274
rect 6773 9222 6783 9274
rect 6783 9222 6829 9274
rect 6533 9220 6589 9222
rect 6613 9220 6669 9222
rect 6693 9220 6749 9222
rect 6773 9220 6829 9222
rect 4302 8186 4358 8188
rect 4382 8186 4438 8188
rect 4462 8186 4518 8188
rect 4542 8186 4598 8188
rect 4302 8134 4348 8186
rect 4348 8134 4358 8186
rect 4382 8134 4412 8186
rect 4412 8134 4424 8186
rect 4424 8134 4438 8186
rect 4462 8134 4476 8186
rect 4476 8134 4488 8186
rect 4488 8134 4518 8186
rect 4542 8134 4552 8186
rect 4552 8134 4598 8186
rect 4302 8132 4358 8134
rect 4382 8132 4438 8134
rect 4462 8132 4518 8134
rect 4542 8132 4598 8134
rect 6533 8186 6589 8188
rect 6613 8186 6669 8188
rect 6693 8186 6749 8188
rect 6773 8186 6829 8188
rect 6533 8134 6579 8186
rect 6579 8134 6589 8186
rect 6613 8134 6643 8186
rect 6643 8134 6655 8186
rect 6655 8134 6669 8186
rect 6693 8134 6707 8186
rect 6707 8134 6719 8186
rect 6719 8134 6749 8186
rect 6773 8134 6783 8186
rect 6783 8134 6829 8186
rect 6533 8132 6589 8134
rect 6613 8132 6669 8134
rect 6693 8132 6749 8134
rect 6773 8132 6829 8134
rect 2731 6554 2787 6556
rect 2811 6554 2867 6556
rect 2891 6554 2947 6556
rect 2971 6554 3027 6556
rect 2731 6502 2777 6554
rect 2777 6502 2787 6554
rect 2811 6502 2841 6554
rect 2841 6502 2853 6554
rect 2853 6502 2867 6554
rect 2891 6502 2905 6554
rect 2905 6502 2917 6554
rect 2917 6502 2947 6554
rect 2971 6502 2981 6554
rect 2981 6502 3027 6554
rect 2731 6500 2787 6502
rect 2811 6500 2867 6502
rect 2891 6500 2947 6502
rect 2971 6500 3027 6502
rect 3606 6332 3608 6352
rect 3608 6332 3660 6352
rect 3660 6332 3662 6352
rect 3606 6296 3662 6332
rect 938 6160 994 6216
rect 2071 6010 2127 6012
rect 2151 6010 2207 6012
rect 2231 6010 2287 6012
rect 2311 6010 2367 6012
rect 2071 5958 2117 6010
rect 2117 5958 2127 6010
rect 2151 5958 2181 6010
rect 2181 5958 2193 6010
rect 2193 5958 2207 6010
rect 2231 5958 2245 6010
rect 2245 5958 2257 6010
rect 2257 5958 2287 6010
rect 2311 5958 2321 6010
rect 2321 5958 2367 6010
rect 2071 5956 2127 5958
rect 2151 5956 2207 5958
rect 2231 5956 2287 5958
rect 2311 5956 2367 5958
rect 4962 7642 5018 7644
rect 5042 7642 5098 7644
rect 5122 7642 5178 7644
rect 5202 7642 5258 7644
rect 4962 7590 5008 7642
rect 5008 7590 5018 7642
rect 5042 7590 5072 7642
rect 5072 7590 5084 7642
rect 5084 7590 5098 7642
rect 5122 7590 5136 7642
rect 5136 7590 5148 7642
rect 5148 7590 5178 7642
rect 5202 7590 5212 7642
rect 5212 7590 5258 7642
rect 4962 7588 5018 7590
rect 5042 7588 5098 7590
rect 5122 7588 5178 7590
rect 5202 7588 5258 7590
rect 4302 7098 4358 7100
rect 4382 7098 4438 7100
rect 4462 7098 4518 7100
rect 4542 7098 4598 7100
rect 4302 7046 4348 7098
rect 4348 7046 4358 7098
rect 4382 7046 4412 7098
rect 4412 7046 4424 7098
rect 4424 7046 4438 7098
rect 4462 7046 4476 7098
rect 4476 7046 4488 7098
rect 4488 7046 4518 7098
rect 4542 7046 4552 7098
rect 4552 7046 4598 7098
rect 4302 7044 4358 7046
rect 4382 7044 4438 7046
rect 4462 7044 4518 7046
rect 4542 7044 4598 7046
rect 2731 5466 2787 5468
rect 2811 5466 2867 5468
rect 2891 5466 2947 5468
rect 2971 5466 3027 5468
rect 2731 5414 2777 5466
rect 2777 5414 2787 5466
rect 2811 5414 2841 5466
rect 2841 5414 2853 5466
rect 2853 5414 2867 5466
rect 2891 5414 2905 5466
rect 2905 5414 2917 5466
rect 2917 5414 2947 5466
rect 2971 5414 2981 5466
rect 2981 5414 3027 5466
rect 2731 5412 2787 5414
rect 2811 5412 2867 5414
rect 2891 5412 2947 5414
rect 2971 5412 3027 5414
rect 1858 4936 1914 4992
rect 2071 4922 2127 4924
rect 2151 4922 2207 4924
rect 2231 4922 2287 4924
rect 2311 4922 2367 4924
rect 2071 4870 2117 4922
rect 2117 4870 2127 4922
rect 2151 4870 2181 4922
rect 2181 4870 2193 4922
rect 2193 4870 2207 4922
rect 2231 4870 2245 4922
rect 2245 4870 2257 4922
rect 2257 4870 2287 4922
rect 2311 4870 2321 4922
rect 2321 4870 2367 4922
rect 2071 4868 2127 4870
rect 2151 4868 2207 4870
rect 2231 4868 2287 4870
rect 2311 4868 2367 4870
rect 2731 4378 2787 4380
rect 2811 4378 2867 4380
rect 2891 4378 2947 4380
rect 2971 4378 3027 4380
rect 2731 4326 2777 4378
rect 2777 4326 2787 4378
rect 2811 4326 2841 4378
rect 2841 4326 2853 4378
rect 2853 4326 2867 4378
rect 2891 4326 2905 4378
rect 2905 4326 2917 4378
rect 2917 4326 2947 4378
rect 2971 4326 2981 4378
rect 2981 4326 3027 4378
rect 2731 4324 2787 4326
rect 2811 4324 2867 4326
rect 2891 4324 2947 4326
rect 2971 4324 3027 4326
rect 2071 3834 2127 3836
rect 2151 3834 2207 3836
rect 2231 3834 2287 3836
rect 2311 3834 2367 3836
rect 2071 3782 2117 3834
rect 2117 3782 2127 3834
rect 2151 3782 2181 3834
rect 2181 3782 2193 3834
rect 2193 3782 2207 3834
rect 2231 3782 2245 3834
rect 2245 3782 2257 3834
rect 2257 3782 2287 3834
rect 2311 3782 2321 3834
rect 2321 3782 2367 3834
rect 2071 3780 2127 3782
rect 2151 3780 2207 3782
rect 2231 3780 2287 3782
rect 2311 3780 2367 3782
rect 2071 2746 2127 2748
rect 2151 2746 2207 2748
rect 2231 2746 2287 2748
rect 2311 2746 2367 2748
rect 2071 2694 2117 2746
rect 2117 2694 2127 2746
rect 2151 2694 2181 2746
rect 2181 2694 2193 2746
rect 2193 2694 2207 2746
rect 2231 2694 2245 2746
rect 2245 2694 2257 2746
rect 2257 2694 2287 2746
rect 2311 2694 2321 2746
rect 2321 2694 2367 2746
rect 2071 2692 2127 2694
rect 2151 2692 2207 2694
rect 2231 2692 2287 2694
rect 2311 2692 2367 2694
rect 4526 6316 4582 6352
rect 4526 6296 4528 6316
rect 4528 6296 4580 6316
rect 4580 6296 4582 6316
rect 4302 6010 4358 6012
rect 4382 6010 4438 6012
rect 4462 6010 4518 6012
rect 4542 6010 4598 6012
rect 4302 5958 4348 6010
rect 4348 5958 4358 6010
rect 4382 5958 4412 6010
rect 4412 5958 4424 6010
rect 4424 5958 4438 6010
rect 4462 5958 4476 6010
rect 4476 5958 4488 6010
rect 4488 5958 4518 6010
rect 4542 5958 4552 6010
rect 4552 5958 4598 6010
rect 4302 5956 4358 5958
rect 4382 5956 4438 5958
rect 4462 5956 4518 5958
rect 4542 5956 4598 5958
rect 4158 5616 4214 5672
rect 4302 4922 4358 4924
rect 4382 4922 4438 4924
rect 4462 4922 4518 4924
rect 4542 4922 4598 4924
rect 4302 4870 4348 4922
rect 4348 4870 4358 4922
rect 4382 4870 4412 4922
rect 4412 4870 4424 4922
rect 4424 4870 4438 4922
rect 4462 4870 4476 4922
rect 4476 4870 4488 4922
rect 4488 4870 4518 4922
rect 4542 4870 4552 4922
rect 4552 4870 4598 4922
rect 4302 4868 4358 4870
rect 4382 4868 4438 4870
rect 4462 4868 4518 4870
rect 4542 4868 4598 4870
rect 2731 3290 2787 3292
rect 2811 3290 2867 3292
rect 2891 3290 2947 3292
rect 2971 3290 3027 3292
rect 2731 3238 2777 3290
rect 2777 3238 2787 3290
rect 2811 3238 2841 3290
rect 2841 3238 2853 3290
rect 2853 3238 2867 3290
rect 2891 3238 2905 3290
rect 2905 3238 2917 3290
rect 2917 3238 2947 3290
rect 2971 3238 2981 3290
rect 2981 3238 3027 3290
rect 2731 3236 2787 3238
rect 2811 3236 2867 3238
rect 2891 3236 2947 3238
rect 2971 3236 3027 3238
rect 4302 3834 4358 3836
rect 4382 3834 4438 3836
rect 4462 3834 4518 3836
rect 4542 3834 4598 3836
rect 4302 3782 4348 3834
rect 4348 3782 4358 3834
rect 4382 3782 4412 3834
rect 4412 3782 4424 3834
rect 4424 3782 4438 3834
rect 4462 3782 4476 3834
rect 4476 3782 4488 3834
rect 4488 3782 4518 3834
rect 4542 3782 4552 3834
rect 4552 3782 4598 3834
rect 4302 3780 4358 3782
rect 4382 3780 4438 3782
rect 4462 3780 4518 3782
rect 4542 3780 4598 3782
rect 4962 6554 5018 6556
rect 5042 6554 5098 6556
rect 5122 6554 5178 6556
rect 5202 6554 5258 6556
rect 4962 6502 5008 6554
rect 5008 6502 5018 6554
rect 5042 6502 5072 6554
rect 5072 6502 5084 6554
rect 5084 6502 5098 6554
rect 5122 6502 5136 6554
rect 5136 6502 5148 6554
rect 5148 6502 5178 6554
rect 5202 6502 5212 6554
rect 5212 6502 5258 6554
rect 4962 6500 5018 6502
rect 5042 6500 5098 6502
rect 5122 6500 5178 6502
rect 5202 6500 5258 6502
rect 4962 5466 5018 5468
rect 5042 5466 5098 5468
rect 5122 5466 5178 5468
rect 5202 5466 5258 5468
rect 4962 5414 5008 5466
rect 5008 5414 5018 5466
rect 5042 5414 5072 5466
rect 5072 5414 5084 5466
rect 5084 5414 5098 5466
rect 5122 5414 5136 5466
rect 5136 5414 5148 5466
rect 5148 5414 5178 5466
rect 5202 5414 5212 5466
rect 5212 5414 5258 5466
rect 4962 5412 5018 5414
rect 5042 5412 5098 5414
rect 5122 5412 5178 5414
rect 5202 5412 5258 5414
rect 4962 4378 5018 4380
rect 5042 4378 5098 4380
rect 5122 4378 5178 4380
rect 5202 4378 5258 4380
rect 4962 4326 5008 4378
rect 5008 4326 5018 4378
rect 5042 4326 5072 4378
rect 5072 4326 5084 4378
rect 5084 4326 5098 4378
rect 5122 4326 5136 4378
rect 5136 4326 5148 4378
rect 5148 4326 5178 4378
rect 5202 4326 5212 4378
rect 5212 4326 5258 4378
rect 4962 4324 5018 4326
rect 5042 4324 5098 4326
rect 5122 4324 5178 4326
rect 5202 4324 5258 4326
rect 4962 3290 5018 3292
rect 5042 3290 5098 3292
rect 5122 3290 5178 3292
rect 5202 3290 5258 3292
rect 4962 3238 5008 3290
rect 5008 3238 5018 3290
rect 5042 3238 5072 3290
rect 5072 3238 5084 3290
rect 5084 3238 5098 3290
rect 5122 3238 5136 3290
rect 5136 3238 5148 3290
rect 5148 3238 5178 3290
rect 5202 3238 5212 3290
rect 5212 3238 5258 3290
rect 4962 3236 5018 3238
rect 5042 3236 5098 3238
rect 5122 3236 5178 3238
rect 5202 3236 5258 3238
rect 4302 2746 4358 2748
rect 4382 2746 4438 2748
rect 4462 2746 4518 2748
rect 4542 2746 4598 2748
rect 4302 2694 4348 2746
rect 4348 2694 4358 2746
rect 4382 2694 4412 2746
rect 4412 2694 4424 2746
rect 4424 2694 4438 2746
rect 4462 2694 4476 2746
rect 4476 2694 4488 2746
rect 4488 2694 4518 2746
rect 4542 2694 4552 2746
rect 4552 2694 4598 2746
rect 4302 2692 4358 2694
rect 4382 2692 4438 2694
rect 4462 2692 4518 2694
rect 4542 2692 4598 2694
rect 1490 1536 1546 1592
rect 2731 2202 2787 2204
rect 2811 2202 2867 2204
rect 2891 2202 2947 2204
rect 2971 2202 3027 2204
rect 2731 2150 2777 2202
rect 2777 2150 2787 2202
rect 2811 2150 2841 2202
rect 2841 2150 2853 2202
rect 2853 2150 2867 2202
rect 2891 2150 2905 2202
rect 2905 2150 2917 2202
rect 2917 2150 2947 2202
rect 2971 2150 2981 2202
rect 2981 2150 3027 2202
rect 2731 2148 2787 2150
rect 2811 2148 2867 2150
rect 2891 2148 2947 2150
rect 2971 2148 3027 2150
rect 7193 8730 7249 8732
rect 7273 8730 7329 8732
rect 7353 8730 7409 8732
rect 7433 8730 7489 8732
rect 7193 8678 7239 8730
rect 7239 8678 7249 8730
rect 7273 8678 7303 8730
rect 7303 8678 7315 8730
rect 7315 8678 7329 8730
rect 7353 8678 7367 8730
rect 7367 8678 7379 8730
rect 7379 8678 7409 8730
rect 7433 8678 7443 8730
rect 7443 8678 7489 8730
rect 7193 8676 7249 8678
rect 7273 8676 7329 8678
rect 7353 8676 7409 8678
rect 7433 8676 7489 8678
rect 7193 7642 7249 7644
rect 7273 7642 7329 7644
rect 7353 7642 7409 7644
rect 7433 7642 7489 7644
rect 7193 7590 7239 7642
rect 7239 7590 7249 7642
rect 7273 7590 7303 7642
rect 7303 7590 7315 7642
rect 7315 7590 7329 7642
rect 7353 7590 7367 7642
rect 7367 7590 7379 7642
rect 7379 7590 7409 7642
rect 7433 7590 7443 7642
rect 7443 7590 7489 7642
rect 7193 7588 7249 7590
rect 7273 7588 7329 7590
rect 7353 7588 7409 7590
rect 7433 7588 7489 7590
rect 6533 7098 6589 7100
rect 6613 7098 6669 7100
rect 6693 7098 6749 7100
rect 6773 7098 6829 7100
rect 6533 7046 6579 7098
rect 6579 7046 6589 7098
rect 6613 7046 6643 7098
rect 6643 7046 6655 7098
rect 6655 7046 6669 7098
rect 6693 7046 6707 7098
rect 6707 7046 6719 7098
rect 6719 7046 6749 7098
rect 6773 7046 6783 7098
rect 6783 7046 6829 7098
rect 6533 7044 6589 7046
rect 6613 7044 6669 7046
rect 6693 7044 6749 7046
rect 6773 7044 6829 7046
rect 6533 6010 6589 6012
rect 6613 6010 6669 6012
rect 6693 6010 6749 6012
rect 6773 6010 6829 6012
rect 6533 5958 6579 6010
rect 6579 5958 6589 6010
rect 6613 5958 6643 6010
rect 6643 5958 6655 6010
rect 6655 5958 6669 6010
rect 6693 5958 6707 6010
rect 6707 5958 6719 6010
rect 6719 5958 6749 6010
rect 6773 5958 6783 6010
rect 6783 5958 6829 6010
rect 6533 5956 6589 5958
rect 6613 5956 6669 5958
rect 6693 5956 6749 5958
rect 6773 5956 6829 5958
rect 6533 4922 6589 4924
rect 6613 4922 6669 4924
rect 6693 4922 6749 4924
rect 6773 4922 6829 4924
rect 6533 4870 6579 4922
rect 6579 4870 6589 4922
rect 6613 4870 6643 4922
rect 6643 4870 6655 4922
rect 6655 4870 6669 4922
rect 6693 4870 6707 4922
rect 6707 4870 6719 4922
rect 6719 4870 6749 4922
rect 6773 4870 6783 4922
rect 6783 4870 6829 4922
rect 6533 4868 6589 4870
rect 6613 4868 6669 4870
rect 6693 4868 6749 4870
rect 6773 4868 6829 4870
rect 9402 12280 9458 12336
rect 9424 10906 9480 10908
rect 9504 10906 9560 10908
rect 9584 10906 9640 10908
rect 9664 10906 9720 10908
rect 9424 10854 9470 10906
rect 9470 10854 9480 10906
rect 9504 10854 9534 10906
rect 9534 10854 9546 10906
rect 9546 10854 9560 10906
rect 9584 10854 9598 10906
rect 9598 10854 9610 10906
rect 9610 10854 9640 10906
rect 9664 10854 9674 10906
rect 9674 10854 9720 10906
rect 9424 10852 9480 10854
rect 9504 10852 9560 10854
rect 9584 10852 9640 10854
rect 9664 10852 9720 10854
rect 8764 10362 8820 10364
rect 8844 10362 8900 10364
rect 8924 10362 8980 10364
rect 9004 10362 9060 10364
rect 8764 10310 8810 10362
rect 8810 10310 8820 10362
rect 8844 10310 8874 10362
rect 8874 10310 8886 10362
rect 8886 10310 8900 10362
rect 8924 10310 8938 10362
rect 8938 10310 8950 10362
rect 8950 10310 8980 10362
rect 9004 10310 9014 10362
rect 9014 10310 9060 10362
rect 8764 10308 8820 10310
rect 8844 10308 8900 10310
rect 8924 10308 8980 10310
rect 9004 10308 9060 10310
rect 8764 9274 8820 9276
rect 8844 9274 8900 9276
rect 8924 9274 8980 9276
rect 9004 9274 9060 9276
rect 8764 9222 8810 9274
rect 8810 9222 8820 9274
rect 8844 9222 8874 9274
rect 8874 9222 8886 9274
rect 8886 9222 8900 9274
rect 8924 9222 8938 9274
rect 8938 9222 8950 9274
rect 8950 9222 8980 9274
rect 9004 9222 9014 9274
rect 9014 9222 9060 9274
rect 8764 9220 8820 9222
rect 8844 9220 8900 9222
rect 8924 9220 8980 9222
rect 9004 9220 9060 9222
rect 7193 6554 7249 6556
rect 7273 6554 7329 6556
rect 7353 6554 7409 6556
rect 7433 6554 7489 6556
rect 7193 6502 7239 6554
rect 7239 6502 7249 6554
rect 7273 6502 7303 6554
rect 7303 6502 7315 6554
rect 7315 6502 7329 6554
rect 7353 6502 7367 6554
rect 7367 6502 7379 6554
rect 7379 6502 7409 6554
rect 7433 6502 7443 6554
rect 7443 6502 7489 6554
rect 7193 6500 7249 6502
rect 7273 6500 7329 6502
rect 7353 6500 7409 6502
rect 7433 6500 7489 6502
rect 7193 5466 7249 5468
rect 7273 5466 7329 5468
rect 7353 5466 7409 5468
rect 7433 5466 7489 5468
rect 7193 5414 7239 5466
rect 7239 5414 7249 5466
rect 7273 5414 7303 5466
rect 7303 5414 7315 5466
rect 7315 5414 7329 5466
rect 7353 5414 7367 5466
rect 7367 5414 7379 5466
rect 7379 5414 7409 5466
rect 7433 5414 7443 5466
rect 7443 5414 7489 5466
rect 7193 5412 7249 5414
rect 7273 5412 7329 5414
rect 7353 5412 7409 5414
rect 7433 5412 7489 5414
rect 6533 3834 6589 3836
rect 6613 3834 6669 3836
rect 6693 3834 6749 3836
rect 6773 3834 6829 3836
rect 6533 3782 6579 3834
rect 6579 3782 6589 3834
rect 6613 3782 6643 3834
rect 6643 3782 6655 3834
rect 6655 3782 6669 3834
rect 6693 3782 6707 3834
rect 6707 3782 6719 3834
rect 6719 3782 6749 3834
rect 6773 3782 6783 3834
rect 6783 3782 6829 3834
rect 6533 3780 6589 3782
rect 6613 3780 6669 3782
rect 6693 3780 6749 3782
rect 6773 3780 6829 3782
rect 7193 4378 7249 4380
rect 7273 4378 7329 4380
rect 7353 4378 7409 4380
rect 7433 4378 7489 4380
rect 7193 4326 7239 4378
rect 7239 4326 7249 4378
rect 7273 4326 7303 4378
rect 7303 4326 7315 4378
rect 7315 4326 7329 4378
rect 7353 4326 7367 4378
rect 7367 4326 7379 4378
rect 7379 4326 7409 4378
rect 7433 4326 7443 4378
rect 7443 4326 7489 4378
rect 7193 4324 7249 4326
rect 7273 4324 7329 4326
rect 7353 4324 7409 4326
rect 7433 4324 7489 4326
rect 7193 3290 7249 3292
rect 7273 3290 7329 3292
rect 7353 3290 7409 3292
rect 7433 3290 7489 3292
rect 7193 3238 7239 3290
rect 7239 3238 7249 3290
rect 7273 3238 7303 3290
rect 7303 3238 7315 3290
rect 7315 3238 7329 3290
rect 7353 3238 7367 3290
rect 7367 3238 7379 3290
rect 7379 3238 7409 3290
rect 7433 3238 7443 3290
rect 7443 3238 7489 3290
rect 7193 3236 7249 3238
rect 7273 3236 7329 3238
rect 7353 3236 7409 3238
rect 7433 3236 7489 3238
rect 9424 9818 9480 9820
rect 9504 9818 9560 9820
rect 9584 9818 9640 9820
rect 9664 9818 9720 9820
rect 9424 9766 9470 9818
rect 9470 9766 9480 9818
rect 9504 9766 9534 9818
rect 9534 9766 9546 9818
rect 9546 9766 9560 9818
rect 9584 9766 9598 9818
rect 9598 9766 9610 9818
rect 9610 9766 9640 9818
rect 9664 9766 9674 9818
rect 9674 9766 9720 9818
rect 9424 9764 9480 9766
rect 9504 9764 9560 9766
rect 9584 9764 9640 9766
rect 9664 9764 9720 9766
rect 9678 8900 9734 8936
rect 9678 8880 9680 8900
rect 9680 8880 9732 8900
rect 9732 8880 9734 8900
rect 9424 8730 9480 8732
rect 9504 8730 9560 8732
rect 9584 8730 9640 8732
rect 9664 8730 9720 8732
rect 9424 8678 9470 8730
rect 9470 8678 9480 8730
rect 9504 8678 9534 8730
rect 9534 8678 9546 8730
rect 9546 8678 9560 8730
rect 9584 8678 9598 8730
rect 9598 8678 9610 8730
rect 9610 8678 9640 8730
rect 9664 8678 9674 8730
rect 9674 8678 9720 8730
rect 9424 8676 9480 8678
rect 9504 8676 9560 8678
rect 9584 8676 9640 8678
rect 9664 8676 9720 8678
rect 8764 8186 8820 8188
rect 8844 8186 8900 8188
rect 8924 8186 8980 8188
rect 9004 8186 9060 8188
rect 8764 8134 8810 8186
rect 8810 8134 8820 8186
rect 8844 8134 8874 8186
rect 8874 8134 8886 8186
rect 8886 8134 8900 8186
rect 8924 8134 8938 8186
rect 8938 8134 8950 8186
rect 8950 8134 8980 8186
rect 9004 8134 9014 8186
rect 9014 8134 9060 8186
rect 8764 8132 8820 8134
rect 8844 8132 8900 8134
rect 8924 8132 8980 8134
rect 9004 8132 9060 8134
rect 8764 7098 8820 7100
rect 8844 7098 8900 7100
rect 8924 7098 8980 7100
rect 9004 7098 9060 7100
rect 8764 7046 8810 7098
rect 8810 7046 8820 7098
rect 8844 7046 8874 7098
rect 8874 7046 8886 7098
rect 8886 7046 8900 7098
rect 8924 7046 8938 7098
rect 8938 7046 8950 7098
rect 8950 7046 8980 7098
rect 9004 7046 9014 7098
rect 9014 7046 9060 7098
rect 8764 7044 8820 7046
rect 8844 7044 8900 7046
rect 8924 7044 8980 7046
rect 9004 7044 9060 7046
rect 9424 7642 9480 7644
rect 9504 7642 9560 7644
rect 9584 7642 9640 7644
rect 9664 7642 9720 7644
rect 9424 7590 9470 7642
rect 9470 7590 9480 7642
rect 9504 7590 9534 7642
rect 9534 7590 9546 7642
rect 9546 7590 9560 7642
rect 9584 7590 9598 7642
rect 9598 7590 9610 7642
rect 9610 7590 9640 7642
rect 9664 7590 9674 7642
rect 9674 7590 9720 7642
rect 9424 7588 9480 7590
rect 9504 7588 9560 7590
rect 9584 7588 9640 7590
rect 9664 7588 9720 7590
rect 9954 7520 10010 7576
rect 9424 6554 9480 6556
rect 9504 6554 9560 6556
rect 9584 6554 9640 6556
rect 9664 6554 9720 6556
rect 9424 6502 9470 6554
rect 9470 6502 9480 6554
rect 9504 6502 9534 6554
rect 9534 6502 9546 6554
rect 9546 6502 9560 6554
rect 9584 6502 9598 6554
rect 9598 6502 9610 6554
rect 9610 6502 9640 6554
rect 9664 6502 9674 6554
rect 9674 6502 9720 6554
rect 9424 6500 9480 6502
rect 9504 6500 9560 6502
rect 9584 6500 9640 6502
rect 9664 6500 9720 6502
rect 8764 6010 8820 6012
rect 8844 6010 8900 6012
rect 8924 6010 8980 6012
rect 9004 6010 9060 6012
rect 8764 5958 8810 6010
rect 8810 5958 8820 6010
rect 8844 5958 8874 6010
rect 8874 5958 8886 6010
rect 8886 5958 8900 6010
rect 8924 5958 8938 6010
rect 8938 5958 8950 6010
rect 8950 5958 8980 6010
rect 9004 5958 9014 6010
rect 9014 5958 9060 6010
rect 8764 5956 8820 5958
rect 8844 5956 8900 5958
rect 8924 5956 8980 5958
rect 9004 5956 9060 5958
rect 10046 5480 10102 5536
rect 9424 5466 9480 5468
rect 9504 5466 9560 5468
rect 9584 5466 9640 5468
rect 9664 5466 9720 5468
rect 9424 5414 9470 5466
rect 9470 5414 9480 5466
rect 9504 5414 9534 5466
rect 9534 5414 9546 5466
rect 9546 5414 9560 5466
rect 9584 5414 9598 5466
rect 9598 5414 9610 5466
rect 9610 5414 9640 5466
rect 9664 5414 9674 5466
rect 9674 5414 9720 5466
rect 9424 5412 9480 5414
rect 9504 5412 9560 5414
rect 9584 5412 9640 5414
rect 9664 5412 9720 5414
rect 8764 4922 8820 4924
rect 8844 4922 8900 4924
rect 8924 4922 8980 4924
rect 9004 4922 9060 4924
rect 8764 4870 8810 4922
rect 8810 4870 8820 4922
rect 8844 4870 8874 4922
rect 8874 4870 8886 4922
rect 8886 4870 8900 4922
rect 8924 4870 8938 4922
rect 8938 4870 8950 4922
rect 8950 4870 8980 4922
rect 9004 4870 9014 4922
rect 9014 4870 9060 4922
rect 8764 4868 8820 4870
rect 8844 4868 8900 4870
rect 8924 4868 8980 4870
rect 9004 4868 9060 4870
rect 8764 3834 8820 3836
rect 8844 3834 8900 3836
rect 8924 3834 8980 3836
rect 9004 3834 9060 3836
rect 8764 3782 8810 3834
rect 8810 3782 8820 3834
rect 8844 3782 8874 3834
rect 8874 3782 8886 3834
rect 8886 3782 8900 3834
rect 8924 3782 8938 3834
rect 8938 3782 8950 3834
rect 8950 3782 8980 3834
rect 9004 3782 9014 3834
rect 9014 3782 9060 3834
rect 8764 3780 8820 3782
rect 8844 3780 8900 3782
rect 8924 3780 8980 3782
rect 9004 3780 9060 3782
rect 6533 2746 6589 2748
rect 6613 2746 6669 2748
rect 6693 2746 6749 2748
rect 6773 2746 6829 2748
rect 6533 2694 6579 2746
rect 6579 2694 6589 2746
rect 6613 2694 6643 2746
rect 6643 2694 6655 2746
rect 6655 2694 6669 2746
rect 6693 2694 6707 2746
rect 6707 2694 6719 2746
rect 6719 2694 6749 2746
rect 6773 2694 6783 2746
rect 6783 2694 6829 2746
rect 6533 2692 6589 2694
rect 6613 2692 6669 2694
rect 6693 2692 6749 2694
rect 6773 2692 6829 2694
rect 4962 2202 5018 2204
rect 5042 2202 5098 2204
rect 5122 2202 5178 2204
rect 5202 2202 5258 2204
rect 4962 2150 5008 2202
rect 5008 2150 5018 2202
rect 5042 2150 5072 2202
rect 5072 2150 5084 2202
rect 5084 2150 5098 2202
rect 5122 2150 5136 2202
rect 5136 2150 5148 2202
rect 5148 2150 5178 2202
rect 5202 2150 5212 2202
rect 5212 2150 5258 2202
rect 4962 2148 5018 2150
rect 5042 2148 5098 2150
rect 5122 2148 5178 2150
rect 5202 2148 5258 2150
rect 7193 2202 7249 2204
rect 7273 2202 7329 2204
rect 7353 2202 7409 2204
rect 7433 2202 7489 2204
rect 7193 2150 7239 2202
rect 7239 2150 7249 2202
rect 7273 2150 7303 2202
rect 7303 2150 7315 2202
rect 7315 2150 7329 2202
rect 7353 2150 7367 2202
rect 7367 2150 7379 2202
rect 7379 2150 7409 2202
rect 7433 2150 7443 2202
rect 7443 2150 7489 2202
rect 7193 2148 7249 2150
rect 7273 2148 7329 2150
rect 7353 2148 7409 2150
rect 7433 2148 7489 2150
rect 8764 2746 8820 2748
rect 8844 2746 8900 2748
rect 8924 2746 8980 2748
rect 9004 2746 9060 2748
rect 8764 2694 8810 2746
rect 8810 2694 8820 2746
rect 8844 2694 8874 2746
rect 8874 2694 8886 2746
rect 8886 2694 8900 2746
rect 8924 2694 8938 2746
rect 8938 2694 8950 2746
rect 8950 2694 8980 2746
rect 9004 2694 9014 2746
rect 9014 2694 9060 2746
rect 8764 2692 8820 2694
rect 8844 2692 8900 2694
rect 8924 2692 8980 2694
rect 9004 2692 9060 2694
rect 9424 4378 9480 4380
rect 9504 4378 9560 4380
rect 9584 4378 9640 4380
rect 9664 4378 9720 4380
rect 9424 4326 9470 4378
rect 9470 4326 9480 4378
rect 9504 4326 9534 4378
rect 9534 4326 9546 4378
rect 9546 4326 9560 4378
rect 9584 4326 9598 4378
rect 9598 4326 9610 4378
rect 9610 4326 9640 4378
rect 9664 4326 9674 4378
rect 9674 4326 9720 4378
rect 9424 4324 9480 4326
rect 9504 4324 9560 4326
rect 9584 4324 9640 4326
rect 9664 4324 9720 4326
rect 9862 4120 9918 4176
rect 9424 3290 9480 3292
rect 9504 3290 9560 3292
rect 9584 3290 9640 3292
rect 9664 3290 9720 3292
rect 9424 3238 9470 3290
rect 9470 3238 9480 3290
rect 9504 3238 9534 3290
rect 9534 3238 9546 3290
rect 9546 3238 9560 3290
rect 9584 3238 9598 3290
rect 9598 3238 9610 3290
rect 9610 3238 9640 3290
rect 9664 3238 9674 3290
rect 9674 3238 9720 3290
rect 9424 3236 9480 3238
rect 9504 3236 9560 3238
rect 9584 3236 9640 3238
rect 9664 3236 9720 3238
rect 9770 2796 9772 2816
rect 9772 2796 9824 2816
rect 9824 2796 9826 2816
rect 9770 2760 9826 2796
rect 9424 2202 9480 2204
rect 9504 2202 9560 2204
rect 9584 2202 9640 2204
rect 9664 2202 9720 2204
rect 9424 2150 9470 2202
rect 9470 2150 9480 2202
rect 9504 2150 9534 2202
rect 9534 2150 9546 2202
rect 9546 2150 9560 2202
rect 9584 2150 9598 2202
rect 9598 2150 9610 2202
rect 9610 2150 9640 2202
rect 9664 2150 9674 2202
rect 9674 2150 9720 2202
rect 9424 2148 9480 2150
rect 9504 2148 9560 2150
rect 9584 2148 9640 2150
rect 9664 2148 9720 2150
rect 8666 720 8722 776
<< metal3 >>
rect 0 13018 800 13048
rect 3049 13018 3115 13021
rect 0 13016 3115 13018
rect 0 12960 3054 13016
rect 3110 12960 3115 13016
rect 0 12958 3115 12960
rect 0 12928 800 12958
rect 3049 12955 3115 12958
rect 9397 12338 9463 12341
rect 10390 12338 11190 12368
rect 9397 12336 11190 12338
rect 9397 12280 9402 12336
rect 9458 12280 11190 12336
rect 9397 12278 11190 12280
rect 9397 12275 9463 12278
rect 10390 12248 11190 12278
rect 0 11658 800 11688
rect 1577 11658 1643 11661
rect 0 11656 1643 11658
rect 0 11600 1582 11656
rect 1638 11600 1643 11656
rect 0 11598 1643 11600
rect 0 11568 800 11598
rect 1577 11595 1643 11598
rect 10390 10978 11190 11008
rect 9814 10918 11190 10978
rect 2721 10912 3037 10913
rect 2721 10848 2727 10912
rect 2791 10848 2807 10912
rect 2871 10848 2887 10912
rect 2951 10848 2967 10912
rect 3031 10848 3037 10912
rect 2721 10847 3037 10848
rect 4952 10912 5268 10913
rect 4952 10848 4958 10912
rect 5022 10848 5038 10912
rect 5102 10848 5118 10912
rect 5182 10848 5198 10912
rect 5262 10848 5268 10912
rect 4952 10847 5268 10848
rect 7183 10912 7499 10913
rect 7183 10848 7189 10912
rect 7253 10848 7269 10912
rect 7333 10848 7349 10912
rect 7413 10848 7429 10912
rect 7493 10848 7499 10912
rect 7183 10847 7499 10848
rect 9414 10912 9730 10913
rect 9414 10848 9420 10912
rect 9484 10848 9500 10912
rect 9564 10848 9580 10912
rect 9644 10848 9660 10912
rect 9724 10848 9730 10912
rect 9414 10847 9730 10848
rect 8201 10706 8267 10709
rect 9814 10706 9874 10918
rect 10390 10888 11190 10918
rect 8201 10704 9874 10706
rect 8201 10648 8206 10704
rect 8262 10648 9874 10704
rect 8201 10646 9874 10648
rect 8201 10643 8267 10646
rect 2061 10368 2377 10369
rect 2061 10304 2067 10368
rect 2131 10304 2147 10368
rect 2211 10304 2227 10368
rect 2291 10304 2307 10368
rect 2371 10304 2377 10368
rect 2061 10303 2377 10304
rect 4292 10368 4608 10369
rect 4292 10304 4298 10368
rect 4362 10304 4378 10368
rect 4442 10304 4458 10368
rect 4522 10304 4538 10368
rect 4602 10304 4608 10368
rect 4292 10303 4608 10304
rect 6523 10368 6839 10369
rect 6523 10304 6529 10368
rect 6593 10304 6609 10368
rect 6673 10304 6689 10368
rect 6753 10304 6769 10368
rect 6833 10304 6839 10368
rect 6523 10303 6839 10304
rect 8754 10368 9070 10369
rect 8754 10304 8760 10368
rect 8824 10304 8840 10368
rect 8904 10304 8920 10368
rect 8984 10304 9000 10368
rect 9064 10304 9070 10368
rect 8754 10303 9070 10304
rect 2721 9824 3037 9825
rect 2721 9760 2727 9824
rect 2791 9760 2807 9824
rect 2871 9760 2887 9824
rect 2951 9760 2967 9824
rect 3031 9760 3037 9824
rect 2721 9759 3037 9760
rect 4952 9824 5268 9825
rect 4952 9760 4958 9824
rect 5022 9760 5038 9824
rect 5102 9760 5118 9824
rect 5182 9760 5198 9824
rect 5262 9760 5268 9824
rect 4952 9759 5268 9760
rect 7183 9824 7499 9825
rect 7183 9760 7189 9824
rect 7253 9760 7269 9824
rect 7333 9760 7349 9824
rect 7413 9760 7429 9824
rect 7493 9760 7499 9824
rect 7183 9759 7499 9760
rect 9414 9824 9730 9825
rect 9414 9760 9420 9824
rect 9484 9760 9500 9824
rect 9564 9760 9580 9824
rect 9644 9760 9660 9824
rect 9724 9760 9730 9824
rect 9414 9759 9730 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 2061 9280 2377 9281
rect 2061 9216 2067 9280
rect 2131 9216 2147 9280
rect 2211 9216 2227 9280
rect 2291 9216 2307 9280
rect 2371 9216 2377 9280
rect 2061 9215 2377 9216
rect 4292 9280 4608 9281
rect 4292 9216 4298 9280
rect 4362 9216 4378 9280
rect 4442 9216 4458 9280
rect 4522 9216 4538 9280
rect 4602 9216 4608 9280
rect 4292 9215 4608 9216
rect 6523 9280 6839 9281
rect 6523 9216 6529 9280
rect 6593 9216 6609 9280
rect 6673 9216 6689 9280
rect 6753 9216 6769 9280
rect 6833 9216 6839 9280
rect 6523 9215 6839 9216
rect 8754 9280 9070 9281
rect 8754 9216 8760 9280
rect 8824 9216 8840 9280
rect 8904 9216 8920 9280
rect 8984 9216 9000 9280
rect 9064 9216 9070 9280
rect 8754 9215 9070 9216
rect 9673 8938 9739 8941
rect 10390 8938 11190 8968
rect 9673 8936 11190 8938
rect 9673 8880 9678 8936
rect 9734 8880 11190 8936
rect 9673 8878 11190 8880
rect 9673 8875 9739 8878
rect 10390 8848 11190 8878
rect 2721 8736 3037 8737
rect 2721 8672 2727 8736
rect 2791 8672 2807 8736
rect 2871 8672 2887 8736
rect 2951 8672 2967 8736
rect 3031 8672 3037 8736
rect 2721 8671 3037 8672
rect 4952 8736 5268 8737
rect 4952 8672 4958 8736
rect 5022 8672 5038 8736
rect 5102 8672 5118 8736
rect 5182 8672 5198 8736
rect 5262 8672 5268 8736
rect 4952 8671 5268 8672
rect 7183 8736 7499 8737
rect 7183 8672 7189 8736
rect 7253 8672 7269 8736
rect 7333 8672 7349 8736
rect 7413 8672 7429 8736
rect 7493 8672 7499 8736
rect 7183 8671 7499 8672
rect 9414 8736 9730 8737
rect 9414 8672 9420 8736
rect 9484 8672 9500 8736
rect 9564 8672 9580 8736
rect 9644 8672 9660 8736
rect 9724 8672 9730 8736
rect 9414 8671 9730 8672
rect 0 8258 800 8288
rect 933 8258 999 8261
rect 0 8256 999 8258
rect 0 8200 938 8256
rect 994 8200 999 8256
rect 0 8198 999 8200
rect 0 8168 800 8198
rect 933 8195 999 8198
rect 2061 8192 2377 8193
rect 2061 8128 2067 8192
rect 2131 8128 2147 8192
rect 2211 8128 2227 8192
rect 2291 8128 2307 8192
rect 2371 8128 2377 8192
rect 2061 8127 2377 8128
rect 4292 8192 4608 8193
rect 4292 8128 4298 8192
rect 4362 8128 4378 8192
rect 4442 8128 4458 8192
rect 4522 8128 4538 8192
rect 4602 8128 4608 8192
rect 4292 8127 4608 8128
rect 6523 8192 6839 8193
rect 6523 8128 6529 8192
rect 6593 8128 6609 8192
rect 6673 8128 6689 8192
rect 6753 8128 6769 8192
rect 6833 8128 6839 8192
rect 6523 8127 6839 8128
rect 8754 8192 9070 8193
rect 8754 8128 8760 8192
rect 8824 8128 8840 8192
rect 8904 8128 8920 8192
rect 8984 8128 9000 8192
rect 9064 8128 9070 8192
rect 8754 8127 9070 8128
rect 2721 7648 3037 7649
rect 2721 7584 2727 7648
rect 2791 7584 2807 7648
rect 2871 7584 2887 7648
rect 2951 7584 2967 7648
rect 3031 7584 3037 7648
rect 2721 7583 3037 7584
rect 4952 7648 5268 7649
rect 4952 7584 4958 7648
rect 5022 7584 5038 7648
rect 5102 7584 5118 7648
rect 5182 7584 5198 7648
rect 5262 7584 5268 7648
rect 4952 7583 5268 7584
rect 7183 7648 7499 7649
rect 7183 7584 7189 7648
rect 7253 7584 7269 7648
rect 7333 7584 7349 7648
rect 7413 7584 7429 7648
rect 7493 7584 7499 7648
rect 7183 7583 7499 7584
rect 9414 7648 9730 7649
rect 9414 7584 9420 7648
rect 9484 7584 9500 7648
rect 9564 7584 9580 7648
rect 9644 7584 9660 7648
rect 9724 7584 9730 7648
rect 9414 7583 9730 7584
rect 9949 7578 10015 7581
rect 10390 7578 11190 7608
rect 9949 7576 11190 7578
rect 9949 7520 9954 7576
rect 10010 7520 11190 7576
rect 9949 7518 11190 7520
rect 9949 7515 10015 7518
rect 10390 7488 11190 7518
rect 2061 7104 2377 7105
rect 2061 7040 2067 7104
rect 2131 7040 2147 7104
rect 2211 7040 2227 7104
rect 2291 7040 2307 7104
rect 2371 7040 2377 7104
rect 2061 7039 2377 7040
rect 4292 7104 4608 7105
rect 4292 7040 4298 7104
rect 4362 7040 4378 7104
rect 4442 7040 4458 7104
rect 4522 7040 4538 7104
rect 4602 7040 4608 7104
rect 4292 7039 4608 7040
rect 6523 7104 6839 7105
rect 6523 7040 6529 7104
rect 6593 7040 6609 7104
rect 6673 7040 6689 7104
rect 6753 7040 6769 7104
rect 6833 7040 6839 7104
rect 6523 7039 6839 7040
rect 8754 7104 9070 7105
rect 8754 7040 8760 7104
rect 8824 7040 8840 7104
rect 8904 7040 8920 7104
rect 8984 7040 9000 7104
rect 9064 7040 9070 7104
rect 8754 7039 9070 7040
rect 2721 6560 3037 6561
rect 2721 6496 2727 6560
rect 2791 6496 2807 6560
rect 2871 6496 2887 6560
rect 2951 6496 2967 6560
rect 3031 6496 3037 6560
rect 2721 6495 3037 6496
rect 4952 6560 5268 6561
rect 4952 6496 4958 6560
rect 5022 6496 5038 6560
rect 5102 6496 5118 6560
rect 5182 6496 5198 6560
rect 5262 6496 5268 6560
rect 4952 6495 5268 6496
rect 7183 6560 7499 6561
rect 7183 6496 7189 6560
rect 7253 6496 7269 6560
rect 7333 6496 7349 6560
rect 7413 6496 7429 6560
rect 7493 6496 7499 6560
rect 7183 6495 7499 6496
rect 9414 6560 9730 6561
rect 9414 6496 9420 6560
rect 9484 6496 9500 6560
rect 9564 6496 9580 6560
rect 9644 6496 9660 6560
rect 9724 6496 9730 6560
rect 9414 6495 9730 6496
rect 3601 6354 3667 6357
rect 4521 6354 4587 6357
rect 3601 6352 4587 6354
rect 3601 6296 3606 6352
rect 3662 6296 4526 6352
rect 4582 6296 4587 6352
rect 3601 6294 4587 6296
rect 3601 6291 3667 6294
rect 4521 6291 4587 6294
rect 0 6218 800 6248
rect 933 6218 999 6221
rect 0 6216 999 6218
rect 0 6160 938 6216
rect 994 6160 999 6216
rect 0 6158 999 6160
rect 0 6128 800 6158
rect 933 6155 999 6158
rect 2061 6016 2377 6017
rect 2061 5952 2067 6016
rect 2131 5952 2147 6016
rect 2211 5952 2227 6016
rect 2291 5952 2307 6016
rect 2371 5952 2377 6016
rect 2061 5951 2377 5952
rect 4292 6016 4608 6017
rect 4292 5952 4298 6016
rect 4362 5952 4378 6016
rect 4442 5952 4458 6016
rect 4522 5952 4538 6016
rect 4602 5952 4608 6016
rect 4292 5951 4608 5952
rect 6523 6016 6839 6017
rect 6523 5952 6529 6016
rect 6593 5952 6609 6016
rect 6673 5952 6689 6016
rect 6753 5952 6769 6016
rect 6833 5952 6839 6016
rect 6523 5951 6839 5952
rect 8754 6016 9070 6017
rect 8754 5952 8760 6016
rect 8824 5952 8840 6016
rect 8904 5952 8920 6016
rect 8984 5952 9000 6016
rect 9064 5952 9070 6016
rect 8754 5951 9070 5952
rect 3734 5612 3740 5676
rect 3804 5674 3810 5676
rect 4153 5674 4219 5677
rect 3804 5672 4219 5674
rect 3804 5616 4158 5672
rect 4214 5616 4219 5672
rect 3804 5614 4219 5616
rect 3804 5612 3810 5614
rect 4153 5611 4219 5614
rect 10041 5538 10107 5541
rect 10390 5538 11190 5568
rect 10041 5536 11190 5538
rect 10041 5480 10046 5536
rect 10102 5480 11190 5536
rect 10041 5478 11190 5480
rect 10041 5475 10107 5478
rect 2721 5472 3037 5473
rect 2721 5408 2727 5472
rect 2791 5408 2807 5472
rect 2871 5408 2887 5472
rect 2951 5408 2967 5472
rect 3031 5408 3037 5472
rect 2721 5407 3037 5408
rect 4952 5472 5268 5473
rect 4952 5408 4958 5472
rect 5022 5408 5038 5472
rect 5102 5408 5118 5472
rect 5182 5408 5198 5472
rect 5262 5408 5268 5472
rect 4952 5407 5268 5408
rect 7183 5472 7499 5473
rect 7183 5408 7189 5472
rect 7253 5408 7269 5472
rect 7333 5408 7349 5472
rect 7413 5408 7429 5472
rect 7493 5408 7499 5472
rect 7183 5407 7499 5408
rect 9414 5472 9730 5473
rect 9414 5408 9420 5472
rect 9484 5408 9500 5472
rect 9564 5408 9580 5472
rect 9644 5408 9660 5472
rect 9724 5408 9730 5472
rect 10390 5448 11190 5478
rect 9414 5407 9730 5408
rect 1853 4994 1919 4997
rect 982 4992 1919 4994
rect 982 4936 1858 4992
rect 1914 4936 1919 4992
rect 982 4934 1919 4936
rect 0 4858 800 4888
rect 982 4858 1042 4934
rect 1853 4931 1919 4934
rect 2061 4928 2377 4929
rect 2061 4864 2067 4928
rect 2131 4864 2147 4928
rect 2211 4864 2227 4928
rect 2291 4864 2307 4928
rect 2371 4864 2377 4928
rect 2061 4863 2377 4864
rect 4292 4928 4608 4929
rect 4292 4864 4298 4928
rect 4362 4864 4378 4928
rect 4442 4864 4458 4928
rect 4522 4864 4538 4928
rect 4602 4864 4608 4928
rect 4292 4863 4608 4864
rect 6523 4928 6839 4929
rect 6523 4864 6529 4928
rect 6593 4864 6609 4928
rect 6673 4864 6689 4928
rect 6753 4864 6769 4928
rect 6833 4864 6839 4928
rect 6523 4863 6839 4864
rect 8754 4928 9070 4929
rect 8754 4864 8760 4928
rect 8824 4864 8840 4928
rect 8904 4864 8920 4928
rect 8984 4864 9000 4928
rect 9064 4864 9070 4928
rect 8754 4863 9070 4864
rect 0 4798 1042 4858
rect 0 4768 800 4798
rect 2721 4384 3037 4385
rect 2721 4320 2727 4384
rect 2791 4320 2807 4384
rect 2871 4320 2887 4384
rect 2951 4320 2967 4384
rect 3031 4320 3037 4384
rect 2721 4319 3037 4320
rect 4952 4384 5268 4385
rect 4952 4320 4958 4384
rect 5022 4320 5038 4384
rect 5102 4320 5118 4384
rect 5182 4320 5198 4384
rect 5262 4320 5268 4384
rect 4952 4319 5268 4320
rect 7183 4384 7499 4385
rect 7183 4320 7189 4384
rect 7253 4320 7269 4384
rect 7333 4320 7349 4384
rect 7413 4320 7429 4384
rect 7493 4320 7499 4384
rect 7183 4319 7499 4320
rect 9414 4384 9730 4385
rect 9414 4320 9420 4384
rect 9484 4320 9500 4384
rect 9564 4320 9580 4384
rect 9644 4320 9660 4384
rect 9724 4320 9730 4384
rect 9414 4319 9730 4320
rect 9857 4178 9923 4181
rect 10390 4178 11190 4208
rect 9857 4176 11190 4178
rect 9857 4120 9862 4176
rect 9918 4120 11190 4176
rect 9857 4118 11190 4120
rect 9857 4115 9923 4118
rect 10390 4088 11190 4118
rect 2061 3840 2377 3841
rect 2061 3776 2067 3840
rect 2131 3776 2147 3840
rect 2211 3776 2227 3840
rect 2291 3776 2307 3840
rect 2371 3776 2377 3840
rect 2061 3775 2377 3776
rect 4292 3840 4608 3841
rect 4292 3776 4298 3840
rect 4362 3776 4378 3840
rect 4442 3776 4458 3840
rect 4522 3776 4538 3840
rect 4602 3776 4608 3840
rect 4292 3775 4608 3776
rect 6523 3840 6839 3841
rect 6523 3776 6529 3840
rect 6593 3776 6609 3840
rect 6673 3776 6689 3840
rect 6753 3776 6769 3840
rect 6833 3776 6839 3840
rect 6523 3775 6839 3776
rect 8754 3840 9070 3841
rect 8754 3776 8760 3840
rect 8824 3776 8840 3840
rect 8904 3776 8920 3840
rect 8984 3776 9000 3840
rect 9064 3776 9070 3840
rect 8754 3775 9070 3776
rect 2721 3296 3037 3297
rect 2721 3232 2727 3296
rect 2791 3232 2807 3296
rect 2871 3232 2887 3296
rect 2951 3232 2967 3296
rect 3031 3232 3037 3296
rect 2721 3231 3037 3232
rect 4952 3296 5268 3297
rect 4952 3232 4958 3296
rect 5022 3232 5038 3296
rect 5102 3232 5118 3296
rect 5182 3232 5198 3296
rect 5262 3232 5268 3296
rect 4952 3231 5268 3232
rect 7183 3296 7499 3297
rect 7183 3232 7189 3296
rect 7253 3232 7269 3296
rect 7333 3232 7349 3296
rect 7413 3232 7429 3296
rect 7493 3232 7499 3296
rect 7183 3231 7499 3232
rect 9414 3296 9730 3297
rect 9414 3232 9420 3296
rect 9484 3232 9500 3296
rect 9564 3232 9580 3296
rect 9644 3232 9660 3296
rect 9724 3232 9730 3296
rect 9414 3231 9730 3232
rect 3734 2954 3740 2956
rect 1902 2894 3740 2954
rect 0 2818 800 2848
rect 1902 2818 1962 2894
rect 3734 2892 3740 2894
rect 3804 2892 3810 2956
rect 0 2758 1962 2818
rect 9765 2818 9831 2821
rect 10390 2818 11190 2848
rect 9765 2816 11190 2818
rect 9765 2760 9770 2816
rect 9826 2760 11190 2816
rect 9765 2758 11190 2760
rect 0 2728 800 2758
rect 9765 2755 9831 2758
rect 2061 2752 2377 2753
rect 2061 2688 2067 2752
rect 2131 2688 2147 2752
rect 2211 2688 2227 2752
rect 2291 2688 2307 2752
rect 2371 2688 2377 2752
rect 2061 2687 2377 2688
rect 4292 2752 4608 2753
rect 4292 2688 4298 2752
rect 4362 2688 4378 2752
rect 4442 2688 4458 2752
rect 4522 2688 4538 2752
rect 4602 2688 4608 2752
rect 4292 2687 4608 2688
rect 6523 2752 6839 2753
rect 6523 2688 6529 2752
rect 6593 2688 6609 2752
rect 6673 2688 6689 2752
rect 6753 2688 6769 2752
rect 6833 2688 6839 2752
rect 6523 2687 6839 2688
rect 8754 2752 9070 2753
rect 8754 2688 8760 2752
rect 8824 2688 8840 2752
rect 8904 2688 8920 2752
rect 8984 2688 9000 2752
rect 9064 2688 9070 2752
rect 10390 2728 11190 2758
rect 8754 2687 9070 2688
rect 2721 2208 3037 2209
rect 2721 2144 2727 2208
rect 2791 2144 2807 2208
rect 2871 2144 2887 2208
rect 2951 2144 2967 2208
rect 3031 2144 3037 2208
rect 2721 2143 3037 2144
rect 4952 2208 5268 2209
rect 4952 2144 4958 2208
rect 5022 2144 5038 2208
rect 5102 2144 5118 2208
rect 5182 2144 5198 2208
rect 5262 2144 5268 2208
rect 4952 2143 5268 2144
rect 7183 2208 7499 2209
rect 7183 2144 7189 2208
rect 7253 2144 7269 2208
rect 7333 2144 7349 2208
rect 7413 2144 7429 2208
rect 7493 2144 7499 2208
rect 7183 2143 7499 2144
rect 9414 2208 9730 2209
rect 9414 2144 9420 2208
rect 9484 2144 9500 2208
rect 9564 2144 9580 2208
rect 9644 2144 9660 2208
rect 9724 2144 9730 2208
rect 9414 2143 9730 2144
rect 1485 1594 1551 1597
rect 982 1592 1551 1594
rect 982 1536 1490 1592
rect 1546 1536 1551 1592
rect 982 1534 1551 1536
rect 0 1458 800 1488
rect 982 1458 1042 1534
rect 1485 1531 1551 1534
rect 0 1398 1042 1458
rect 0 1368 800 1398
rect 8661 778 8727 781
rect 10390 778 11190 808
rect 8661 776 11190 778
rect 8661 720 8666 776
rect 8722 720 11190 776
rect 8661 718 11190 720
rect 8661 715 8727 718
rect 10390 688 11190 718
<< via3 >>
rect 2727 10908 2791 10912
rect 2727 10852 2731 10908
rect 2731 10852 2787 10908
rect 2787 10852 2791 10908
rect 2727 10848 2791 10852
rect 2807 10908 2871 10912
rect 2807 10852 2811 10908
rect 2811 10852 2867 10908
rect 2867 10852 2871 10908
rect 2807 10848 2871 10852
rect 2887 10908 2951 10912
rect 2887 10852 2891 10908
rect 2891 10852 2947 10908
rect 2947 10852 2951 10908
rect 2887 10848 2951 10852
rect 2967 10908 3031 10912
rect 2967 10852 2971 10908
rect 2971 10852 3027 10908
rect 3027 10852 3031 10908
rect 2967 10848 3031 10852
rect 4958 10908 5022 10912
rect 4958 10852 4962 10908
rect 4962 10852 5018 10908
rect 5018 10852 5022 10908
rect 4958 10848 5022 10852
rect 5038 10908 5102 10912
rect 5038 10852 5042 10908
rect 5042 10852 5098 10908
rect 5098 10852 5102 10908
rect 5038 10848 5102 10852
rect 5118 10908 5182 10912
rect 5118 10852 5122 10908
rect 5122 10852 5178 10908
rect 5178 10852 5182 10908
rect 5118 10848 5182 10852
rect 5198 10908 5262 10912
rect 5198 10852 5202 10908
rect 5202 10852 5258 10908
rect 5258 10852 5262 10908
rect 5198 10848 5262 10852
rect 7189 10908 7253 10912
rect 7189 10852 7193 10908
rect 7193 10852 7249 10908
rect 7249 10852 7253 10908
rect 7189 10848 7253 10852
rect 7269 10908 7333 10912
rect 7269 10852 7273 10908
rect 7273 10852 7329 10908
rect 7329 10852 7333 10908
rect 7269 10848 7333 10852
rect 7349 10908 7413 10912
rect 7349 10852 7353 10908
rect 7353 10852 7409 10908
rect 7409 10852 7413 10908
rect 7349 10848 7413 10852
rect 7429 10908 7493 10912
rect 7429 10852 7433 10908
rect 7433 10852 7489 10908
rect 7489 10852 7493 10908
rect 7429 10848 7493 10852
rect 9420 10908 9484 10912
rect 9420 10852 9424 10908
rect 9424 10852 9480 10908
rect 9480 10852 9484 10908
rect 9420 10848 9484 10852
rect 9500 10908 9564 10912
rect 9500 10852 9504 10908
rect 9504 10852 9560 10908
rect 9560 10852 9564 10908
rect 9500 10848 9564 10852
rect 9580 10908 9644 10912
rect 9580 10852 9584 10908
rect 9584 10852 9640 10908
rect 9640 10852 9644 10908
rect 9580 10848 9644 10852
rect 9660 10908 9724 10912
rect 9660 10852 9664 10908
rect 9664 10852 9720 10908
rect 9720 10852 9724 10908
rect 9660 10848 9724 10852
rect 2067 10364 2131 10368
rect 2067 10308 2071 10364
rect 2071 10308 2127 10364
rect 2127 10308 2131 10364
rect 2067 10304 2131 10308
rect 2147 10364 2211 10368
rect 2147 10308 2151 10364
rect 2151 10308 2207 10364
rect 2207 10308 2211 10364
rect 2147 10304 2211 10308
rect 2227 10364 2291 10368
rect 2227 10308 2231 10364
rect 2231 10308 2287 10364
rect 2287 10308 2291 10364
rect 2227 10304 2291 10308
rect 2307 10364 2371 10368
rect 2307 10308 2311 10364
rect 2311 10308 2367 10364
rect 2367 10308 2371 10364
rect 2307 10304 2371 10308
rect 4298 10364 4362 10368
rect 4298 10308 4302 10364
rect 4302 10308 4358 10364
rect 4358 10308 4362 10364
rect 4298 10304 4362 10308
rect 4378 10364 4442 10368
rect 4378 10308 4382 10364
rect 4382 10308 4438 10364
rect 4438 10308 4442 10364
rect 4378 10304 4442 10308
rect 4458 10364 4522 10368
rect 4458 10308 4462 10364
rect 4462 10308 4518 10364
rect 4518 10308 4522 10364
rect 4458 10304 4522 10308
rect 4538 10364 4602 10368
rect 4538 10308 4542 10364
rect 4542 10308 4598 10364
rect 4598 10308 4602 10364
rect 4538 10304 4602 10308
rect 6529 10364 6593 10368
rect 6529 10308 6533 10364
rect 6533 10308 6589 10364
rect 6589 10308 6593 10364
rect 6529 10304 6593 10308
rect 6609 10364 6673 10368
rect 6609 10308 6613 10364
rect 6613 10308 6669 10364
rect 6669 10308 6673 10364
rect 6609 10304 6673 10308
rect 6689 10364 6753 10368
rect 6689 10308 6693 10364
rect 6693 10308 6749 10364
rect 6749 10308 6753 10364
rect 6689 10304 6753 10308
rect 6769 10364 6833 10368
rect 6769 10308 6773 10364
rect 6773 10308 6829 10364
rect 6829 10308 6833 10364
rect 6769 10304 6833 10308
rect 8760 10364 8824 10368
rect 8760 10308 8764 10364
rect 8764 10308 8820 10364
rect 8820 10308 8824 10364
rect 8760 10304 8824 10308
rect 8840 10364 8904 10368
rect 8840 10308 8844 10364
rect 8844 10308 8900 10364
rect 8900 10308 8904 10364
rect 8840 10304 8904 10308
rect 8920 10364 8984 10368
rect 8920 10308 8924 10364
rect 8924 10308 8980 10364
rect 8980 10308 8984 10364
rect 8920 10304 8984 10308
rect 9000 10364 9064 10368
rect 9000 10308 9004 10364
rect 9004 10308 9060 10364
rect 9060 10308 9064 10364
rect 9000 10304 9064 10308
rect 2727 9820 2791 9824
rect 2727 9764 2731 9820
rect 2731 9764 2787 9820
rect 2787 9764 2791 9820
rect 2727 9760 2791 9764
rect 2807 9820 2871 9824
rect 2807 9764 2811 9820
rect 2811 9764 2867 9820
rect 2867 9764 2871 9820
rect 2807 9760 2871 9764
rect 2887 9820 2951 9824
rect 2887 9764 2891 9820
rect 2891 9764 2947 9820
rect 2947 9764 2951 9820
rect 2887 9760 2951 9764
rect 2967 9820 3031 9824
rect 2967 9764 2971 9820
rect 2971 9764 3027 9820
rect 3027 9764 3031 9820
rect 2967 9760 3031 9764
rect 4958 9820 5022 9824
rect 4958 9764 4962 9820
rect 4962 9764 5018 9820
rect 5018 9764 5022 9820
rect 4958 9760 5022 9764
rect 5038 9820 5102 9824
rect 5038 9764 5042 9820
rect 5042 9764 5098 9820
rect 5098 9764 5102 9820
rect 5038 9760 5102 9764
rect 5118 9820 5182 9824
rect 5118 9764 5122 9820
rect 5122 9764 5178 9820
rect 5178 9764 5182 9820
rect 5118 9760 5182 9764
rect 5198 9820 5262 9824
rect 5198 9764 5202 9820
rect 5202 9764 5258 9820
rect 5258 9764 5262 9820
rect 5198 9760 5262 9764
rect 7189 9820 7253 9824
rect 7189 9764 7193 9820
rect 7193 9764 7249 9820
rect 7249 9764 7253 9820
rect 7189 9760 7253 9764
rect 7269 9820 7333 9824
rect 7269 9764 7273 9820
rect 7273 9764 7329 9820
rect 7329 9764 7333 9820
rect 7269 9760 7333 9764
rect 7349 9820 7413 9824
rect 7349 9764 7353 9820
rect 7353 9764 7409 9820
rect 7409 9764 7413 9820
rect 7349 9760 7413 9764
rect 7429 9820 7493 9824
rect 7429 9764 7433 9820
rect 7433 9764 7489 9820
rect 7489 9764 7493 9820
rect 7429 9760 7493 9764
rect 9420 9820 9484 9824
rect 9420 9764 9424 9820
rect 9424 9764 9480 9820
rect 9480 9764 9484 9820
rect 9420 9760 9484 9764
rect 9500 9820 9564 9824
rect 9500 9764 9504 9820
rect 9504 9764 9560 9820
rect 9560 9764 9564 9820
rect 9500 9760 9564 9764
rect 9580 9820 9644 9824
rect 9580 9764 9584 9820
rect 9584 9764 9640 9820
rect 9640 9764 9644 9820
rect 9580 9760 9644 9764
rect 9660 9820 9724 9824
rect 9660 9764 9664 9820
rect 9664 9764 9720 9820
rect 9720 9764 9724 9820
rect 9660 9760 9724 9764
rect 2067 9276 2131 9280
rect 2067 9220 2071 9276
rect 2071 9220 2127 9276
rect 2127 9220 2131 9276
rect 2067 9216 2131 9220
rect 2147 9276 2211 9280
rect 2147 9220 2151 9276
rect 2151 9220 2207 9276
rect 2207 9220 2211 9276
rect 2147 9216 2211 9220
rect 2227 9276 2291 9280
rect 2227 9220 2231 9276
rect 2231 9220 2287 9276
rect 2287 9220 2291 9276
rect 2227 9216 2291 9220
rect 2307 9276 2371 9280
rect 2307 9220 2311 9276
rect 2311 9220 2367 9276
rect 2367 9220 2371 9276
rect 2307 9216 2371 9220
rect 4298 9276 4362 9280
rect 4298 9220 4302 9276
rect 4302 9220 4358 9276
rect 4358 9220 4362 9276
rect 4298 9216 4362 9220
rect 4378 9276 4442 9280
rect 4378 9220 4382 9276
rect 4382 9220 4438 9276
rect 4438 9220 4442 9276
rect 4378 9216 4442 9220
rect 4458 9276 4522 9280
rect 4458 9220 4462 9276
rect 4462 9220 4518 9276
rect 4518 9220 4522 9276
rect 4458 9216 4522 9220
rect 4538 9276 4602 9280
rect 4538 9220 4542 9276
rect 4542 9220 4598 9276
rect 4598 9220 4602 9276
rect 4538 9216 4602 9220
rect 6529 9276 6593 9280
rect 6529 9220 6533 9276
rect 6533 9220 6589 9276
rect 6589 9220 6593 9276
rect 6529 9216 6593 9220
rect 6609 9276 6673 9280
rect 6609 9220 6613 9276
rect 6613 9220 6669 9276
rect 6669 9220 6673 9276
rect 6609 9216 6673 9220
rect 6689 9276 6753 9280
rect 6689 9220 6693 9276
rect 6693 9220 6749 9276
rect 6749 9220 6753 9276
rect 6689 9216 6753 9220
rect 6769 9276 6833 9280
rect 6769 9220 6773 9276
rect 6773 9220 6829 9276
rect 6829 9220 6833 9276
rect 6769 9216 6833 9220
rect 8760 9276 8824 9280
rect 8760 9220 8764 9276
rect 8764 9220 8820 9276
rect 8820 9220 8824 9276
rect 8760 9216 8824 9220
rect 8840 9276 8904 9280
rect 8840 9220 8844 9276
rect 8844 9220 8900 9276
rect 8900 9220 8904 9276
rect 8840 9216 8904 9220
rect 8920 9276 8984 9280
rect 8920 9220 8924 9276
rect 8924 9220 8980 9276
rect 8980 9220 8984 9276
rect 8920 9216 8984 9220
rect 9000 9276 9064 9280
rect 9000 9220 9004 9276
rect 9004 9220 9060 9276
rect 9060 9220 9064 9276
rect 9000 9216 9064 9220
rect 2727 8732 2791 8736
rect 2727 8676 2731 8732
rect 2731 8676 2787 8732
rect 2787 8676 2791 8732
rect 2727 8672 2791 8676
rect 2807 8732 2871 8736
rect 2807 8676 2811 8732
rect 2811 8676 2867 8732
rect 2867 8676 2871 8732
rect 2807 8672 2871 8676
rect 2887 8732 2951 8736
rect 2887 8676 2891 8732
rect 2891 8676 2947 8732
rect 2947 8676 2951 8732
rect 2887 8672 2951 8676
rect 2967 8732 3031 8736
rect 2967 8676 2971 8732
rect 2971 8676 3027 8732
rect 3027 8676 3031 8732
rect 2967 8672 3031 8676
rect 4958 8732 5022 8736
rect 4958 8676 4962 8732
rect 4962 8676 5018 8732
rect 5018 8676 5022 8732
rect 4958 8672 5022 8676
rect 5038 8732 5102 8736
rect 5038 8676 5042 8732
rect 5042 8676 5098 8732
rect 5098 8676 5102 8732
rect 5038 8672 5102 8676
rect 5118 8732 5182 8736
rect 5118 8676 5122 8732
rect 5122 8676 5178 8732
rect 5178 8676 5182 8732
rect 5118 8672 5182 8676
rect 5198 8732 5262 8736
rect 5198 8676 5202 8732
rect 5202 8676 5258 8732
rect 5258 8676 5262 8732
rect 5198 8672 5262 8676
rect 7189 8732 7253 8736
rect 7189 8676 7193 8732
rect 7193 8676 7249 8732
rect 7249 8676 7253 8732
rect 7189 8672 7253 8676
rect 7269 8732 7333 8736
rect 7269 8676 7273 8732
rect 7273 8676 7329 8732
rect 7329 8676 7333 8732
rect 7269 8672 7333 8676
rect 7349 8732 7413 8736
rect 7349 8676 7353 8732
rect 7353 8676 7409 8732
rect 7409 8676 7413 8732
rect 7349 8672 7413 8676
rect 7429 8732 7493 8736
rect 7429 8676 7433 8732
rect 7433 8676 7489 8732
rect 7489 8676 7493 8732
rect 7429 8672 7493 8676
rect 9420 8732 9484 8736
rect 9420 8676 9424 8732
rect 9424 8676 9480 8732
rect 9480 8676 9484 8732
rect 9420 8672 9484 8676
rect 9500 8732 9564 8736
rect 9500 8676 9504 8732
rect 9504 8676 9560 8732
rect 9560 8676 9564 8732
rect 9500 8672 9564 8676
rect 9580 8732 9644 8736
rect 9580 8676 9584 8732
rect 9584 8676 9640 8732
rect 9640 8676 9644 8732
rect 9580 8672 9644 8676
rect 9660 8732 9724 8736
rect 9660 8676 9664 8732
rect 9664 8676 9720 8732
rect 9720 8676 9724 8732
rect 9660 8672 9724 8676
rect 2067 8188 2131 8192
rect 2067 8132 2071 8188
rect 2071 8132 2127 8188
rect 2127 8132 2131 8188
rect 2067 8128 2131 8132
rect 2147 8188 2211 8192
rect 2147 8132 2151 8188
rect 2151 8132 2207 8188
rect 2207 8132 2211 8188
rect 2147 8128 2211 8132
rect 2227 8188 2291 8192
rect 2227 8132 2231 8188
rect 2231 8132 2287 8188
rect 2287 8132 2291 8188
rect 2227 8128 2291 8132
rect 2307 8188 2371 8192
rect 2307 8132 2311 8188
rect 2311 8132 2367 8188
rect 2367 8132 2371 8188
rect 2307 8128 2371 8132
rect 4298 8188 4362 8192
rect 4298 8132 4302 8188
rect 4302 8132 4358 8188
rect 4358 8132 4362 8188
rect 4298 8128 4362 8132
rect 4378 8188 4442 8192
rect 4378 8132 4382 8188
rect 4382 8132 4438 8188
rect 4438 8132 4442 8188
rect 4378 8128 4442 8132
rect 4458 8188 4522 8192
rect 4458 8132 4462 8188
rect 4462 8132 4518 8188
rect 4518 8132 4522 8188
rect 4458 8128 4522 8132
rect 4538 8188 4602 8192
rect 4538 8132 4542 8188
rect 4542 8132 4598 8188
rect 4598 8132 4602 8188
rect 4538 8128 4602 8132
rect 6529 8188 6593 8192
rect 6529 8132 6533 8188
rect 6533 8132 6589 8188
rect 6589 8132 6593 8188
rect 6529 8128 6593 8132
rect 6609 8188 6673 8192
rect 6609 8132 6613 8188
rect 6613 8132 6669 8188
rect 6669 8132 6673 8188
rect 6609 8128 6673 8132
rect 6689 8188 6753 8192
rect 6689 8132 6693 8188
rect 6693 8132 6749 8188
rect 6749 8132 6753 8188
rect 6689 8128 6753 8132
rect 6769 8188 6833 8192
rect 6769 8132 6773 8188
rect 6773 8132 6829 8188
rect 6829 8132 6833 8188
rect 6769 8128 6833 8132
rect 8760 8188 8824 8192
rect 8760 8132 8764 8188
rect 8764 8132 8820 8188
rect 8820 8132 8824 8188
rect 8760 8128 8824 8132
rect 8840 8188 8904 8192
rect 8840 8132 8844 8188
rect 8844 8132 8900 8188
rect 8900 8132 8904 8188
rect 8840 8128 8904 8132
rect 8920 8188 8984 8192
rect 8920 8132 8924 8188
rect 8924 8132 8980 8188
rect 8980 8132 8984 8188
rect 8920 8128 8984 8132
rect 9000 8188 9064 8192
rect 9000 8132 9004 8188
rect 9004 8132 9060 8188
rect 9060 8132 9064 8188
rect 9000 8128 9064 8132
rect 2727 7644 2791 7648
rect 2727 7588 2731 7644
rect 2731 7588 2787 7644
rect 2787 7588 2791 7644
rect 2727 7584 2791 7588
rect 2807 7644 2871 7648
rect 2807 7588 2811 7644
rect 2811 7588 2867 7644
rect 2867 7588 2871 7644
rect 2807 7584 2871 7588
rect 2887 7644 2951 7648
rect 2887 7588 2891 7644
rect 2891 7588 2947 7644
rect 2947 7588 2951 7644
rect 2887 7584 2951 7588
rect 2967 7644 3031 7648
rect 2967 7588 2971 7644
rect 2971 7588 3027 7644
rect 3027 7588 3031 7644
rect 2967 7584 3031 7588
rect 4958 7644 5022 7648
rect 4958 7588 4962 7644
rect 4962 7588 5018 7644
rect 5018 7588 5022 7644
rect 4958 7584 5022 7588
rect 5038 7644 5102 7648
rect 5038 7588 5042 7644
rect 5042 7588 5098 7644
rect 5098 7588 5102 7644
rect 5038 7584 5102 7588
rect 5118 7644 5182 7648
rect 5118 7588 5122 7644
rect 5122 7588 5178 7644
rect 5178 7588 5182 7644
rect 5118 7584 5182 7588
rect 5198 7644 5262 7648
rect 5198 7588 5202 7644
rect 5202 7588 5258 7644
rect 5258 7588 5262 7644
rect 5198 7584 5262 7588
rect 7189 7644 7253 7648
rect 7189 7588 7193 7644
rect 7193 7588 7249 7644
rect 7249 7588 7253 7644
rect 7189 7584 7253 7588
rect 7269 7644 7333 7648
rect 7269 7588 7273 7644
rect 7273 7588 7329 7644
rect 7329 7588 7333 7644
rect 7269 7584 7333 7588
rect 7349 7644 7413 7648
rect 7349 7588 7353 7644
rect 7353 7588 7409 7644
rect 7409 7588 7413 7644
rect 7349 7584 7413 7588
rect 7429 7644 7493 7648
rect 7429 7588 7433 7644
rect 7433 7588 7489 7644
rect 7489 7588 7493 7644
rect 7429 7584 7493 7588
rect 9420 7644 9484 7648
rect 9420 7588 9424 7644
rect 9424 7588 9480 7644
rect 9480 7588 9484 7644
rect 9420 7584 9484 7588
rect 9500 7644 9564 7648
rect 9500 7588 9504 7644
rect 9504 7588 9560 7644
rect 9560 7588 9564 7644
rect 9500 7584 9564 7588
rect 9580 7644 9644 7648
rect 9580 7588 9584 7644
rect 9584 7588 9640 7644
rect 9640 7588 9644 7644
rect 9580 7584 9644 7588
rect 9660 7644 9724 7648
rect 9660 7588 9664 7644
rect 9664 7588 9720 7644
rect 9720 7588 9724 7644
rect 9660 7584 9724 7588
rect 2067 7100 2131 7104
rect 2067 7044 2071 7100
rect 2071 7044 2127 7100
rect 2127 7044 2131 7100
rect 2067 7040 2131 7044
rect 2147 7100 2211 7104
rect 2147 7044 2151 7100
rect 2151 7044 2207 7100
rect 2207 7044 2211 7100
rect 2147 7040 2211 7044
rect 2227 7100 2291 7104
rect 2227 7044 2231 7100
rect 2231 7044 2287 7100
rect 2287 7044 2291 7100
rect 2227 7040 2291 7044
rect 2307 7100 2371 7104
rect 2307 7044 2311 7100
rect 2311 7044 2367 7100
rect 2367 7044 2371 7100
rect 2307 7040 2371 7044
rect 4298 7100 4362 7104
rect 4298 7044 4302 7100
rect 4302 7044 4358 7100
rect 4358 7044 4362 7100
rect 4298 7040 4362 7044
rect 4378 7100 4442 7104
rect 4378 7044 4382 7100
rect 4382 7044 4438 7100
rect 4438 7044 4442 7100
rect 4378 7040 4442 7044
rect 4458 7100 4522 7104
rect 4458 7044 4462 7100
rect 4462 7044 4518 7100
rect 4518 7044 4522 7100
rect 4458 7040 4522 7044
rect 4538 7100 4602 7104
rect 4538 7044 4542 7100
rect 4542 7044 4598 7100
rect 4598 7044 4602 7100
rect 4538 7040 4602 7044
rect 6529 7100 6593 7104
rect 6529 7044 6533 7100
rect 6533 7044 6589 7100
rect 6589 7044 6593 7100
rect 6529 7040 6593 7044
rect 6609 7100 6673 7104
rect 6609 7044 6613 7100
rect 6613 7044 6669 7100
rect 6669 7044 6673 7100
rect 6609 7040 6673 7044
rect 6689 7100 6753 7104
rect 6689 7044 6693 7100
rect 6693 7044 6749 7100
rect 6749 7044 6753 7100
rect 6689 7040 6753 7044
rect 6769 7100 6833 7104
rect 6769 7044 6773 7100
rect 6773 7044 6829 7100
rect 6829 7044 6833 7100
rect 6769 7040 6833 7044
rect 8760 7100 8824 7104
rect 8760 7044 8764 7100
rect 8764 7044 8820 7100
rect 8820 7044 8824 7100
rect 8760 7040 8824 7044
rect 8840 7100 8904 7104
rect 8840 7044 8844 7100
rect 8844 7044 8900 7100
rect 8900 7044 8904 7100
rect 8840 7040 8904 7044
rect 8920 7100 8984 7104
rect 8920 7044 8924 7100
rect 8924 7044 8980 7100
rect 8980 7044 8984 7100
rect 8920 7040 8984 7044
rect 9000 7100 9064 7104
rect 9000 7044 9004 7100
rect 9004 7044 9060 7100
rect 9060 7044 9064 7100
rect 9000 7040 9064 7044
rect 2727 6556 2791 6560
rect 2727 6500 2731 6556
rect 2731 6500 2787 6556
rect 2787 6500 2791 6556
rect 2727 6496 2791 6500
rect 2807 6556 2871 6560
rect 2807 6500 2811 6556
rect 2811 6500 2867 6556
rect 2867 6500 2871 6556
rect 2807 6496 2871 6500
rect 2887 6556 2951 6560
rect 2887 6500 2891 6556
rect 2891 6500 2947 6556
rect 2947 6500 2951 6556
rect 2887 6496 2951 6500
rect 2967 6556 3031 6560
rect 2967 6500 2971 6556
rect 2971 6500 3027 6556
rect 3027 6500 3031 6556
rect 2967 6496 3031 6500
rect 4958 6556 5022 6560
rect 4958 6500 4962 6556
rect 4962 6500 5018 6556
rect 5018 6500 5022 6556
rect 4958 6496 5022 6500
rect 5038 6556 5102 6560
rect 5038 6500 5042 6556
rect 5042 6500 5098 6556
rect 5098 6500 5102 6556
rect 5038 6496 5102 6500
rect 5118 6556 5182 6560
rect 5118 6500 5122 6556
rect 5122 6500 5178 6556
rect 5178 6500 5182 6556
rect 5118 6496 5182 6500
rect 5198 6556 5262 6560
rect 5198 6500 5202 6556
rect 5202 6500 5258 6556
rect 5258 6500 5262 6556
rect 5198 6496 5262 6500
rect 7189 6556 7253 6560
rect 7189 6500 7193 6556
rect 7193 6500 7249 6556
rect 7249 6500 7253 6556
rect 7189 6496 7253 6500
rect 7269 6556 7333 6560
rect 7269 6500 7273 6556
rect 7273 6500 7329 6556
rect 7329 6500 7333 6556
rect 7269 6496 7333 6500
rect 7349 6556 7413 6560
rect 7349 6500 7353 6556
rect 7353 6500 7409 6556
rect 7409 6500 7413 6556
rect 7349 6496 7413 6500
rect 7429 6556 7493 6560
rect 7429 6500 7433 6556
rect 7433 6500 7489 6556
rect 7489 6500 7493 6556
rect 7429 6496 7493 6500
rect 9420 6556 9484 6560
rect 9420 6500 9424 6556
rect 9424 6500 9480 6556
rect 9480 6500 9484 6556
rect 9420 6496 9484 6500
rect 9500 6556 9564 6560
rect 9500 6500 9504 6556
rect 9504 6500 9560 6556
rect 9560 6500 9564 6556
rect 9500 6496 9564 6500
rect 9580 6556 9644 6560
rect 9580 6500 9584 6556
rect 9584 6500 9640 6556
rect 9640 6500 9644 6556
rect 9580 6496 9644 6500
rect 9660 6556 9724 6560
rect 9660 6500 9664 6556
rect 9664 6500 9720 6556
rect 9720 6500 9724 6556
rect 9660 6496 9724 6500
rect 2067 6012 2131 6016
rect 2067 5956 2071 6012
rect 2071 5956 2127 6012
rect 2127 5956 2131 6012
rect 2067 5952 2131 5956
rect 2147 6012 2211 6016
rect 2147 5956 2151 6012
rect 2151 5956 2207 6012
rect 2207 5956 2211 6012
rect 2147 5952 2211 5956
rect 2227 6012 2291 6016
rect 2227 5956 2231 6012
rect 2231 5956 2287 6012
rect 2287 5956 2291 6012
rect 2227 5952 2291 5956
rect 2307 6012 2371 6016
rect 2307 5956 2311 6012
rect 2311 5956 2367 6012
rect 2367 5956 2371 6012
rect 2307 5952 2371 5956
rect 4298 6012 4362 6016
rect 4298 5956 4302 6012
rect 4302 5956 4358 6012
rect 4358 5956 4362 6012
rect 4298 5952 4362 5956
rect 4378 6012 4442 6016
rect 4378 5956 4382 6012
rect 4382 5956 4438 6012
rect 4438 5956 4442 6012
rect 4378 5952 4442 5956
rect 4458 6012 4522 6016
rect 4458 5956 4462 6012
rect 4462 5956 4518 6012
rect 4518 5956 4522 6012
rect 4458 5952 4522 5956
rect 4538 6012 4602 6016
rect 4538 5956 4542 6012
rect 4542 5956 4598 6012
rect 4598 5956 4602 6012
rect 4538 5952 4602 5956
rect 6529 6012 6593 6016
rect 6529 5956 6533 6012
rect 6533 5956 6589 6012
rect 6589 5956 6593 6012
rect 6529 5952 6593 5956
rect 6609 6012 6673 6016
rect 6609 5956 6613 6012
rect 6613 5956 6669 6012
rect 6669 5956 6673 6012
rect 6609 5952 6673 5956
rect 6689 6012 6753 6016
rect 6689 5956 6693 6012
rect 6693 5956 6749 6012
rect 6749 5956 6753 6012
rect 6689 5952 6753 5956
rect 6769 6012 6833 6016
rect 6769 5956 6773 6012
rect 6773 5956 6829 6012
rect 6829 5956 6833 6012
rect 6769 5952 6833 5956
rect 8760 6012 8824 6016
rect 8760 5956 8764 6012
rect 8764 5956 8820 6012
rect 8820 5956 8824 6012
rect 8760 5952 8824 5956
rect 8840 6012 8904 6016
rect 8840 5956 8844 6012
rect 8844 5956 8900 6012
rect 8900 5956 8904 6012
rect 8840 5952 8904 5956
rect 8920 6012 8984 6016
rect 8920 5956 8924 6012
rect 8924 5956 8980 6012
rect 8980 5956 8984 6012
rect 8920 5952 8984 5956
rect 9000 6012 9064 6016
rect 9000 5956 9004 6012
rect 9004 5956 9060 6012
rect 9060 5956 9064 6012
rect 9000 5952 9064 5956
rect 3740 5612 3804 5676
rect 2727 5468 2791 5472
rect 2727 5412 2731 5468
rect 2731 5412 2787 5468
rect 2787 5412 2791 5468
rect 2727 5408 2791 5412
rect 2807 5468 2871 5472
rect 2807 5412 2811 5468
rect 2811 5412 2867 5468
rect 2867 5412 2871 5468
rect 2807 5408 2871 5412
rect 2887 5468 2951 5472
rect 2887 5412 2891 5468
rect 2891 5412 2947 5468
rect 2947 5412 2951 5468
rect 2887 5408 2951 5412
rect 2967 5468 3031 5472
rect 2967 5412 2971 5468
rect 2971 5412 3027 5468
rect 3027 5412 3031 5468
rect 2967 5408 3031 5412
rect 4958 5468 5022 5472
rect 4958 5412 4962 5468
rect 4962 5412 5018 5468
rect 5018 5412 5022 5468
rect 4958 5408 5022 5412
rect 5038 5468 5102 5472
rect 5038 5412 5042 5468
rect 5042 5412 5098 5468
rect 5098 5412 5102 5468
rect 5038 5408 5102 5412
rect 5118 5468 5182 5472
rect 5118 5412 5122 5468
rect 5122 5412 5178 5468
rect 5178 5412 5182 5468
rect 5118 5408 5182 5412
rect 5198 5468 5262 5472
rect 5198 5412 5202 5468
rect 5202 5412 5258 5468
rect 5258 5412 5262 5468
rect 5198 5408 5262 5412
rect 7189 5468 7253 5472
rect 7189 5412 7193 5468
rect 7193 5412 7249 5468
rect 7249 5412 7253 5468
rect 7189 5408 7253 5412
rect 7269 5468 7333 5472
rect 7269 5412 7273 5468
rect 7273 5412 7329 5468
rect 7329 5412 7333 5468
rect 7269 5408 7333 5412
rect 7349 5468 7413 5472
rect 7349 5412 7353 5468
rect 7353 5412 7409 5468
rect 7409 5412 7413 5468
rect 7349 5408 7413 5412
rect 7429 5468 7493 5472
rect 7429 5412 7433 5468
rect 7433 5412 7489 5468
rect 7489 5412 7493 5468
rect 7429 5408 7493 5412
rect 9420 5468 9484 5472
rect 9420 5412 9424 5468
rect 9424 5412 9480 5468
rect 9480 5412 9484 5468
rect 9420 5408 9484 5412
rect 9500 5468 9564 5472
rect 9500 5412 9504 5468
rect 9504 5412 9560 5468
rect 9560 5412 9564 5468
rect 9500 5408 9564 5412
rect 9580 5468 9644 5472
rect 9580 5412 9584 5468
rect 9584 5412 9640 5468
rect 9640 5412 9644 5468
rect 9580 5408 9644 5412
rect 9660 5468 9724 5472
rect 9660 5412 9664 5468
rect 9664 5412 9720 5468
rect 9720 5412 9724 5468
rect 9660 5408 9724 5412
rect 2067 4924 2131 4928
rect 2067 4868 2071 4924
rect 2071 4868 2127 4924
rect 2127 4868 2131 4924
rect 2067 4864 2131 4868
rect 2147 4924 2211 4928
rect 2147 4868 2151 4924
rect 2151 4868 2207 4924
rect 2207 4868 2211 4924
rect 2147 4864 2211 4868
rect 2227 4924 2291 4928
rect 2227 4868 2231 4924
rect 2231 4868 2287 4924
rect 2287 4868 2291 4924
rect 2227 4864 2291 4868
rect 2307 4924 2371 4928
rect 2307 4868 2311 4924
rect 2311 4868 2367 4924
rect 2367 4868 2371 4924
rect 2307 4864 2371 4868
rect 4298 4924 4362 4928
rect 4298 4868 4302 4924
rect 4302 4868 4358 4924
rect 4358 4868 4362 4924
rect 4298 4864 4362 4868
rect 4378 4924 4442 4928
rect 4378 4868 4382 4924
rect 4382 4868 4438 4924
rect 4438 4868 4442 4924
rect 4378 4864 4442 4868
rect 4458 4924 4522 4928
rect 4458 4868 4462 4924
rect 4462 4868 4518 4924
rect 4518 4868 4522 4924
rect 4458 4864 4522 4868
rect 4538 4924 4602 4928
rect 4538 4868 4542 4924
rect 4542 4868 4598 4924
rect 4598 4868 4602 4924
rect 4538 4864 4602 4868
rect 6529 4924 6593 4928
rect 6529 4868 6533 4924
rect 6533 4868 6589 4924
rect 6589 4868 6593 4924
rect 6529 4864 6593 4868
rect 6609 4924 6673 4928
rect 6609 4868 6613 4924
rect 6613 4868 6669 4924
rect 6669 4868 6673 4924
rect 6609 4864 6673 4868
rect 6689 4924 6753 4928
rect 6689 4868 6693 4924
rect 6693 4868 6749 4924
rect 6749 4868 6753 4924
rect 6689 4864 6753 4868
rect 6769 4924 6833 4928
rect 6769 4868 6773 4924
rect 6773 4868 6829 4924
rect 6829 4868 6833 4924
rect 6769 4864 6833 4868
rect 8760 4924 8824 4928
rect 8760 4868 8764 4924
rect 8764 4868 8820 4924
rect 8820 4868 8824 4924
rect 8760 4864 8824 4868
rect 8840 4924 8904 4928
rect 8840 4868 8844 4924
rect 8844 4868 8900 4924
rect 8900 4868 8904 4924
rect 8840 4864 8904 4868
rect 8920 4924 8984 4928
rect 8920 4868 8924 4924
rect 8924 4868 8980 4924
rect 8980 4868 8984 4924
rect 8920 4864 8984 4868
rect 9000 4924 9064 4928
rect 9000 4868 9004 4924
rect 9004 4868 9060 4924
rect 9060 4868 9064 4924
rect 9000 4864 9064 4868
rect 2727 4380 2791 4384
rect 2727 4324 2731 4380
rect 2731 4324 2787 4380
rect 2787 4324 2791 4380
rect 2727 4320 2791 4324
rect 2807 4380 2871 4384
rect 2807 4324 2811 4380
rect 2811 4324 2867 4380
rect 2867 4324 2871 4380
rect 2807 4320 2871 4324
rect 2887 4380 2951 4384
rect 2887 4324 2891 4380
rect 2891 4324 2947 4380
rect 2947 4324 2951 4380
rect 2887 4320 2951 4324
rect 2967 4380 3031 4384
rect 2967 4324 2971 4380
rect 2971 4324 3027 4380
rect 3027 4324 3031 4380
rect 2967 4320 3031 4324
rect 4958 4380 5022 4384
rect 4958 4324 4962 4380
rect 4962 4324 5018 4380
rect 5018 4324 5022 4380
rect 4958 4320 5022 4324
rect 5038 4380 5102 4384
rect 5038 4324 5042 4380
rect 5042 4324 5098 4380
rect 5098 4324 5102 4380
rect 5038 4320 5102 4324
rect 5118 4380 5182 4384
rect 5118 4324 5122 4380
rect 5122 4324 5178 4380
rect 5178 4324 5182 4380
rect 5118 4320 5182 4324
rect 5198 4380 5262 4384
rect 5198 4324 5202 4380
rect 5202 4324 5258 4380
rect 5258 4324 5262 4380
rect 5198 4320 5262 4324
rect 7189 4380 7253 4384
rect 7189 4324 7193 4380
rect 7193 4324 7249 4380
rect 7249 4324 7253 4380
rect 7189 4320 7253 4324
rect 7269 4380 7333 4384
rect 7269 4324 7273 4380
rect 7273 4324 7329 4380
rect 7329 4324 7333 4380
rect 7269 4320 7333 4324
rect 7349 4380 7413 4384
rect 7349 4324 7353 4380
rect 7353 4324 7409 4380
rect 7409 4324 7413 4380
rect 7349 4320 7413 4324
rect 7429 4380 7493 4384
rect 7429 4324 7433 4380
rect 7433 4324 7489 4380
rect 7489 4324 7493 4380
rect 7429 4320 7493 4324
rect 9420 4380 9484 4384
rect 9420 4324 9424 4380
rect 9424 4324 9480 4380
rect 9480 4324 9484 4380
rect 9420 4320 9484 4324
rect 9500 4380 9564 4384
rect 9500 4324 9504 4380
rect 9504 4324 9560 4380
rect 9560 4324 9564 4380
rect 9500 4320 9564 4324
rect 9580 4380 9644 4384
rect 9580 4324 9584 4380
rect 9584 4324 9640 4380
rect 9640 4324 9644 4380
rect 9580 4320 9644 4324
rect 9660 4380 9724 4384
rect 9660 4324 9664 4380
rect 9664 4324 9720 4380
rect 9720 4324 9724 4380
rect 9660 4320 9724 4324
rect 2067 3836 2131 3840
rect 2067 3780 2071 3836
rect 2071 3780 2127 3836
rect 2127 3780 2131 3836
rect 2067 3776 2131 3780
rect 2147 3836 2211 3840
rect 2147 3780 2151 3836
rect 2151 3780 2207 3836
rect 2207 3780 2211 3836
rect 2147 3776 2211 3780
rect 2227 3836 2291 3840
rect 2227 3780 2231 3836
rect 2231 3780 2287 3836
rect 2287 3780 2291 3836
rect 2227 3776 2291 3780
rect 2307 3836 2371 3840
rect 2307 3780 2311 3836
rect 2311 3780 2367 3836
rect 2367 3780 2371 3836
rect 2307 3776 2371 3780
rect 4298 3836 4362 3840
rect 4298 3780 4302 3836
rect 4302 3780 4358 3836
rect 4358 3780 4362 3836
rect 4298 3776 4362 3780
rect 4378 3836 4442 3840
rect 4378 3780 4382 3836
rect 4382 3780 4438 3836
rect 4438 3780 4442 3836
rect 4378 3776 4442 3780
rect 4458 3836 4522 3840
rect 4458 3780 4462 3836
rect 4462 3780 4518 3836
rect 4518 3780 4522 3836
rect 4458 3776 4522 3780
rect 4538 3836 4602 3840
rect 4538 3780 4542 3836
rect 4542 3780 4598 3836
rect 4598 3780 4602 3836
rect 4538 3776 4602 3780
rect 6529 3836 6593 3840
rect 6529 3780 6533 3836
rect 6533 3780 6589 3836
rect 6589 3780 6593 3836
rect 6529 3776 6593 3780
rect 6609 3836 6673 3840
rect 6609 3780 6613 3836
rect 6613 3780 6669 3836
rect 6669 3780 6673 3836
rect 6609 3776 6673 3780
rect 6689 3836 6753 3840
rect 6689 3780 6693 3836
rect 6693 3780 6749 3836
rect 6749 3780 6753 3836
rect 6689 3776 6753 3780
rect 6769 3836 6833 3840
rect 6769 3780 6773 3836
rect 6773 3780 6829 3836
rect 6829 3780 6833 3836
rect 6769 3776 6833 3780
rect 8760 3836 8824 3840
rect 8760 3780 8764 3836
rect 8764 3780 8820 3836
rect 8820 3780 8824 3836
rect 8760 3776 8824 3780
rect 8840 3836 8904 3840
rect 8840 3780 8844 3836
rect 8844 3780 8900 3836
rect 8900 3780 8904 3836
rect 8840 3776 8904 3780
rect 8920 3836 8984 3840
rect 8920 3780 8924 3836
rect 8924 3780 8980 3836
rect 8980 3780 8984 3836
rect 8920 3776 8984 3780
rect 9000 3836 9064 3840
rect 9000 3780 9004 3836
rect 9004 3780 9060 3836
rect 9060 3780 9064 3836
rect 9000 3776 9064 3780
rect 2727 3292 2791 3296
rect 2727 3236 2731 3292
rect 2731 3236 2787 3292
rect 2787 3236 2791 3292
rect 2727 3232 2791 3236
rect 2807 3292 2871 3296
rect 2807 3236 2811 3292
rect 2811 3236 2867 3292
rect 2867 3236 2871 3292
rect 2807 3232 2871 3236
rect 2887 3292 2951 3296
rect 2887 3236 2891 3292
rect 2891 3236 2947 3292
rect 2947 3236 2951 3292
rect 2887 3232 2951 3236
rect 2967 3292 3031 3296
rect 2967 3236 2971 3292
rect 2971 3236 3027 3292
rect 3027 3236 3031 3292
rect 2967 3232 3031 3236
rect 4958 3292 5022 3296
rect 4958 3236 4962 3292
rect 4962 3236 5018 3292
rect 5018 3236 5022 3292
rect 4958 3232 5022 3236
rect 5038 3292 5102 3296
rect 5038 3236 5042 3292
rect 5042 3236 5098 3292
rect 5098 3236 5102 3292
rect 5038 3232 5102 3236
rect 5118 3292 5182 3296
rect 5118 3236 5122 3292
rect 5122 3236 5178 3292
rect 5178 3236 5182 3292
rect 5118 3232 5182 3236
rect 5198 3292 5262 3296
rect 5198 3236 5202 3292
rect 5202 3236 5258 3292
rect 5258 3236 5262 3292
rect 5198 3232 5262 3236
rect 7189 3292 7253 3296
rect 7189 3236 7193 3292
rect 7193 3236 7249 3292
rect 7249 3236 7253 3292
rect 7189 3232 7253 3236
rect 7269 3292 7333 3296
rect 7269 3236 7273 3292
rect 7273 3236 7329 3292
rect 7329 3236 7333 3292
rect 7269 3232 7333 3236
rect 7349 3292 7413 3296
rect 7349 3236 7353 3292
rect 7353 3236 7409 3292
rect 7409 3236 7413 3292
rect 7349 3232 7413 3236
rect 7429 3292 7493 3296
rect 7429 3236 7433 3292
rect 7433 3236 7489 3292
rect 7489 3236 7493 3292
rect 7429 3232 7493 3236
rect 9420 3292 9484 3296
rect 9420 3236 9424 3292
rect 9424 3236 9480 3292
rect 9480 3236 9484 3292
rect 9420 3232 9484 3236
rect 9500 3292 9564 3296
rect 9500 3236 9504 3292
rect 9504 3236 9560 3292
rect 9560 3236 9564 3292
rect 9500 3232 9564 3236
rect 9580 3292 9644 3296
rect 9580 3236 9584 3292
rect 9584 3236 9640 3292
rect 9640 3236 9644 3292
rect 9580 3232 9644 3236
rect 9660 3292 9724 3296
rect 9660 3236 9664 3292
rect 9664 3236 9720 3292
rect 9720 3236 9724 3292
rect 9660 3232 9724 3236
rect 3740 2892 3804 2956
rect 2067 2748 2131 2752
rect 2067 2692 2071 2748
rect 2071 2692 2127 2748
rect 2127 2692 2131 2748
rect 2067 2688 2131 2692
rect 2147 2748 2211 2752
rect 2147 2692 2151 2748
rect 2151 2692 2207 2748
rect 2207 2692 2211 2748
rect 2147 2688 2211 2692
rect 2227 2748 2291 2752
rect 2227 2692 2231 2748
rect 2231 2692 2287 2748
rect 2287 2692 2291 2748
rect 2227 2688 2291 2692
rect 2307 2748 2371 2752
rect 2307 2692 2311 2748
rect 2311 2692 2367 2748
rect 2367 2692 2371 2748
rect 2307 2688 2371 2692
rect 4298 2748 4362 2752
rect 4298 2692 4302 2748
rect 4302 2692 4358 2748
rect 4358 2692 4362 2748
rect 4298 2688 4362 2692
rect 4378 2748 4442 2752
rect 4378 2692 4382 2748
rect 4382 2692 4438 2748
rect 4438 2692 4442 2748
rect 4378 2688 4442 2692
rect 4458 2748 4522 2752
rect 4458 2692 4462 2748
rect 4462 2692 4518 2748
rect 4518 2692 4522 2748
rect 4458 2688 4522 2692
rect 4538 2748 4602 2752
rect 4538 2692 4542 2748
rect 4542 2692 4598 2748
rect 4598 2692 4602 2748
rect 4538 2688 4602 2692
rect 6529 2748 6593 2752
rect 6529 2692 6533 2748
rect 6533 2692 6589 2748
rect 6589 2692 6593 2748
rect 6529 2688 6593 2692
rect 6609 2748 6673 2752
rect 6609 2692 6613 2748
rect 6613 2692 6669 2748
rect 6669 2692 6673 2748
rect 6609 2688 6673 2692
rect 6689 2748 6753 2752
rect 6689 2692 6693 2748
rect 6693 2692 6749 2748
rect 6749 2692 6753 2748
rect 6689 2688 6753 2692
rect 6769 2748 6833 2752
rect 6769 2692 6773 2748
rect 6773 2692 6829 2748
rect 6829 2692 6833 2748
rect 6769 2688 6833 2692
rect 8760 2748 8824 2752
rect 8760 2692 8764 2748
rect 8764 2692 8820 2748
rect 8820 2692 8824 2748
rect 8760 2688 8824 2692
rect 8840 2748 8904 2752
rect 8840 2692 8844 2748
rect 8844 2692 8900 2748
rect 8900 2692 8904 2748
rect 8840 2688 8904 2692
rect 8920 2748 8984 2752
rect 8920 2692 8924 2748
rect 8924 2692 8980 2748
rect 8980 2692 8984 2748
rect 8920 2688 8984 2692
rect 9000 2748 9064 2752
rect 9000 2692 9004 2748
rect 9004 2692 9060 2748
rect 9060 2692 9064 2748
rect 9000 2688 9064 2692
rect 2727 2204 2791 2208
rect 2727 2148 2731 2204
rect 2731 2148 2787 2204
rect 2787 2148 2791 2204
rect 2727 2144 2791 2148
rect 2807 2204 2871 2208
rect 2807 2148 2811 2204
rect 2811 2148 2867 2204
rect 2867 2148 2871 2204
rect 2807 2144 2871 2148
rect 2887 2204 2951 2208
rect 2887 2148 2891 2204
rect 2891 2148 2947 2204
rect 2947 2148 2951 2204
rect 2887 2144 2951 2148
rect 2967 2204 3031 2208
rect 2967 2148 2971 2204
rect 2971 2148 3027 2204
rect 3027 2148 3031 2204
rect 2967 2144 3031 2148
rect 4958 2204 5022 2208
rect 4958 2148 4962 2204
rect 4962 2148 5018 2204
rect 5018 2148 5022 2204
rect 4958 2144 5022 2148
rect 5038 2204 5102 2208
rect 5038 2148 5042 2204
rect 5042 2148 5098 2204
rect 5098 2148 5102 2204
rect 5038 2144 5102 2148
rect 5118 2204 5182 2208
rect 5118 2148 5122 2204
rect 5122 2148 5178 2204
rect 5178 2148 5182 2204
rect 5118 2144 5182 2148
rect 5198 2204 5262 2208
rect 5198 2148 5202 2204
rect 5202 2148 5258 2204
rect 5258 2148 5262 2204
rect 5198 2144 5262 2148
rect 7189 2204 7253 2208
rect 7189 2148 7193 2204
rect 7193 2148 7249 2204
rect 7249 2148 7253 2204
rect 7189 2144 7253 2148
rect 7269 2204 7333 2208
rect 7269 2148 7273 2204
rect 7273 2148 7329 2204
rect 7329 2148 7333 2204
rect 7269 2144 7333 2148
rect 7349 2204 7413 2208
rect 7349 2148 7353 2204
rect 7353 2148 7409 2204
rect 7409 2148 7413 2204
rect 7349 2144 7413 2148
rect 7429 2204 7493 2208
rect 7429 2148 7433 2204
rect 7433 2148 7489 2204
rect 7489 2148 7493 2204
rect 7429 2144 7493 2148
rect 9420 2204 9484 2208
rect 9420 2148 9424 2204
rect 9424 2148 9480 2204
rect 9480 2148 9484 2204
rect 9420 2144 9484 2148
rect 9500 2204 9564 2208
rect 9500 2148 9504 2204
rect 9504 2148 9560 2204
rect 9560 2148 9564 2204
rect 9500 2144 9564 2148
rect 9580 2204 9644 2208
rect 9580 2148 9584 2204
rect 9584 2148 9640 2204
rect 9640 2148 9644 2204
rect 9580 2144 9644 2148
rect 9660 2204 9724 2208
rect 9660 2148 9664 2204
rect 9664 2148 9720 2204
rect 9720 2148 9724 2204
rect 9660 2144 9724 2148
<< metal4 >>
rect 2059 10368 2379 10928
rect 2059 10304 2067 10368
rect 2131 10304 2147 10368
rect 2211 10304 2227 10368
rect 2291 10304 2307 10368
rect 2371 10304 2379 10368
rect 2059 9906 2379 10304
rect 2059 9670 2101 9906
rect 2337 9670 2379 9906
rect 2059 9280 2379 9670
rect 2059 9216 2067 9280
rect 2131 9216 2147 9280
rect 2211 9216 2227 9280
rect 2291 9216 2307 9280
rect 2371 9216 2379 9280
rect 2059 8192 2379 9216
rect 2059 8128 2067 8192
rect 2131 8128 2147 8192
rect 2211 8128 2227 8192
rect 2291 8128 2307 8192
rect 2371 8128 2379 8192
rect 2059 7731 2379 8128
rect 2059 7495 2101 7731
rect 2337 7495 2379 7731
rect 2059 7104 2379 7495
rect 2059 7040 2067 7104
rect 2131 7040 2147 7104
rect 2211 7040 2227 7104
rect 2291 7040 2307 7104
rect 2371 7040 2379 7104
rect 2059 6016 2379 7040
rect 2059 5952 2067 6016
rect 2131 5952 2147 6016
rect 2211 5952 2227 6016
rect 2291 5952 2307 6016
rect 2371 5952 2379 6016
rect 2059 5556 2379 5952
rect 2059 5320 2101 5556
rect 2337 5320 2379 5556
rect 2059 4928 2379 5320
rect 2059 4864 2067 4928
rect 2131 4864 2147 4928
rect 2211 4864 2227 4928
rect 2291 4864 2307 4928
rect 2371 4864 2379 4928
rect 2059 3840 2379 4864
rect 2059 3776 2067 3840
rect 2131 3776 2147 3840
rect 2211 3776 2227 3840
rect 2291 3776 2307 3840
rect 2371 3776 2379 3840
rect 2059 3381 2379 3776
rect 2059 3145 2101 3381
rect 2337 3145 2379 3381
rect 2059 2752 2379 3145
rect 2059 2688 2067 2752
rect 2131 2688 2147 2752
rect 2211 2688 2227 2752
rect 2291 2688 2307 2752
rect 2371 2688 2379 2752
rect 2059 2128 2379 2688
rect 2719 10912 3039 10928
rect 2719 10848 2727 10912
rect 2791 10848 2807 10912
rect 2871 10848 2887 10912
rect 2951 10848 2967 10912
rect 3031 10848 3039 10912
rect 2719 10566 3039 10848
rect 2719 10330 2761 10566
rect 2997 10330 3039 10566
rect 2719 9824 3039 10330
rect 2719 9760 2727 9824
rect 2791 9760 2807 9824
rect 2871 9760 2887 9824
rect 2951 9760 2967 9824
rect 3031 9760 3039 9824
rect 2719 8736 3039 9760
rect 2719 8672 2727 8736
rect 2791 8672 2807 8736
rect 2871 8672 2887 8736
rect 2951 8672 2967 8736
rect 3031 8672 3039 8736
rect 2719 8391 3039 8672
rect 2719 8155 2761 8391
rect 2997 8155 3039 8391
rect 2719 7648 3039 8155
rect 2719 7584 2727 7648
rect 2791 7584 2807 7648
rect 2871 7584 2887 7648
rect 2951 7584 2967 7648
rect 3031 7584 3039 7648
rect 2719 6560 3039 7584
rect 2719 6496 2727 6560
rect 2791 6496 2807 6560
rect 2871 6496 2887 6560
rect 2951 6496 2967 6560
rect 3031 6496 3039 6560
rect 2719 6216 3039 6496
rect 2719 5980 2761 6216
rect 2997 5980 3039 6216
rect 2719 5472 3039 5980
rect 4290 10368 4610 10928
rect 4290 10304 4298 10368
rect 4362 10304 4378 10368
rect 4442 10304 4458 10368
rect 4522 10304 4538 10368
rect 4602 10304 4610 10368
rect 4290 9906 4610 10304
rect 4290 9670 4332 9906
rect 4568 9670 4610 9906
rect 4290 9280 4610 9670
rect 4290 9216 4298 9280
rect 4362 9216 4378 9280
rect 4442 9216 4458 9280
rect 4522 9216 4538 9280
rect 4602 9216 4610 9280
rect 4290 8192 4610 9216
rect 4290 8128 4298 8192
rect 4362 8128 4378 8192
rect 4442 8128 4458 8192
rect 4522 8128 4538 8192
rect 4602 8128 4610 8192
rect 4290 7731 4610 8128
rect 4290 7495 4332 7731
rect 4568 7495 4610 7731
rect 4290 7104 4610 7495
rect 4290 7040 4298 7104
rect 4362 7040 4378 7104
rect 4442 7040 4458 7104
rect 4522 7040 4538 7104
rect 4602 7040 4610 7104
rect 4290 6016 4610 7040
rect 4290 5952 4298 6016
rect 4362 5952 4378 6016
rect 4442 5952 4458 6016
rect 4522 5952 4538 6016
rect 4602 5952 4610 6016
rect 3739 5676 3805 5677
rect 3739 5612 3740 5676
rect 3804 5612 3805 5676
rect 3739 5611 3805 5612
rect 2719 5408 2727 5472
rect 2791 5408 2807 5472
rect 2871 5408 2887 5472
rect 2951 5408 2967 5472
rect 3031 5408 3039 5472
rect 2719 4384 3039 5408
rect 2719 4320 2727 4384
rect 2791 4320 2807 4384
rect 2871 4320 2887 4384
rect 2951 4320 2967 4384
rect 3031 4320 3039 4384
rect 2719 4041 3039 4320
rect 2719 3805 2761 4041
rect 2997 3805 3039 4041
rect 2719 3296 3039 3805
rect 2719 3232 2727 3296
rect 2791 3232 2807 3296
rect 2871 3232 2887 3296
rect 2951 3232 2967 3296
rect 3031 3232 3039 3296
rect 2719 2208 3039 3232
rect 3742 2957 3802 5611
rect 4290 5556 4610 5952
rect 4290 5320 4332 5556
rect 4568 5320 4610 5556
rect 4290 4928 4610 5320
rect 4290 4864 4298 4928
rect 4362 4864 4378 4928
rect 4442 4864 4458 4928
rect 4522 4864 4538 4928
rect 4602 4864 4610 4928
rect 4290 3840 4610 4864
rect 4290 3776 4298 3840
rect 4362 3776 4378 3840
rect 4442 3776 4458 3840
rect 4522 3776 4538 3840
rect 4602 3776 4610 3840
rect 4290 3381 4610 3776
rect 4290 3145 4332 3381
rect 4568 3145 4610 3381
rect 3739 2956 3805 2957
rect 3739 2892 3740 2956
rect 3804 2892 3805 2956
rect 3739 2891 3805 2892
rect 2719 2144 2727 2208
rect 2791 2144 2807 2208
rect 2871 2144 2887 2208
rect 2951 2144 2967 2208
rect 3031 2144 3039 2208
rect 2719 2128 3039 2144
rect 4290 2752 4610 3145
rect 4290 2688 4298 2752
rect 4362 2688 4378 2752
rect 4442 2688 4458 2752
rect 4522 2688 4538 2752
rect 4602 2688 4610 2752
rect 4290 2128 4610 2688
rect 4950 10912 5270 10928
rect 4950 10848 4958 10912
rect 5022 10848 5038 10912
rect 5102 10848 5118 10912
rect 5182 10848 5198 10912
rect 5262 10848 5270 10912
rect 4950 10566 5270 10848
rect 4950 10330 4992 10566
rect 5228 10330 5270 10566
rect 4950 9824 5270 10330
rect 4950 9760 4958 9824
rect 5022 9760 5038 9824
rect 5102 9760 5118 9824
rect 5182 9760 5198 9824
rect 5262 9760 5270 9824
rect 4950 8736 5270 9760
rect 4950 8672 4958 8736
rect 5022 8672 5038 8736
rect 5102 8672 5118 8736
rect 5182 8672 5198 8736
rect 5262 8672 5270 8736
rect 4950 8391 5270 8672
rect 4950 8155 4992 8391
rect 5228 8155 5270 8391
rect 4950 7648 5270 8155
rect 4950 7584 4958 7648
rect 5022 7584 5038 7648
rect 5102 7584 5118 7648
rect 5182 7584 5198 7648
rect 5262 7584 5270 7648
rect 4950 6560 5270 7584
rect 4950 6496 4958 6560
rect 5022 6496 5038 6560
rect 5102 6496 5118 6560
rect 5182 6496 5198 6560
rect 5262 6496 5270 6560
rect 4950 6216 5270 6496
rect 4950 5980 4992 6216
rect 5228 5980 5270 6216
rect 4950 5472 5270 5980
rect 4950 5408 4958 5472
rect 5022 5408 5038 5472
rect 5102 5408 5118 5472
rect 5182 5408 5198 5472
rect 5262 5408 5270 5472
rect 4950 4384 5270 5408
rect 4950 4320 4958 4384
rect 5022 4320 5038 4384
rect 5102 4320 5118 4384
rect 5182 4320 5198 4384
rect 5262 4320 5270 4384
rect 4950 4041 5270 4320
rect 4950 3805 4992 4041
rect 5228 3805 5270 4041
rect 4950 3296 5270 3805
rect 4950 3232 4958 3296
rect 5022 3232 5038 3296
rect 5102 3232 5118 3296
rect 5182 3232 5198 3296
rect 5262 3232 5270 3296
rect 4950 2208 5270 3232
rect 4950 2144 4958 2208
rect 5022 2144 5038 2208
rect 5102 2144 5118 2208
rect 5182 2144 5198 2208
rect 5262 2144 5270 2208
rect 4950 2128 5270 2144
rect 6521 10368 6841 10928
rect 6521 10304 6529 10368
rect 6593 10304 6609 10368
rect 6673 10304 6689 10368
rect 6753 10304 6769 10368
rect 6833 10304 6841 10368
rect 6521 9906 6841 10304
rect 6521 9670 6563 9906
rect 6799 9670 6841 9906
rect 6521 9280 6841 9670
rect 6521 9216 6529 9280
rect 6593 9216 6609 9280
rect 6673 9216 6689 9280
rect 6753 9216 6769 9280
rect 6833 9216 6841 9280
rect 6521 8192 6841 9216
rect 6521 8128 6529 8192
rect 6593 8128 6609 8192
rect 6673 8128 6689 8192
rect 6753 8128 6769 8192
rect 6833 8128 6841 8192
rect 6521 7731 6841 8128
rect 6521 7495 6563 7731
rect 6799 7495 6841 7731
rect 6521 7104 6841 7495
rect 6521 7040 6529 7104
rect 6593 7040 6609 7104
rect 6673 7040 6689 7104
rect 6753 7040 6769 7104
rect 6833 7040 6841 7104
rect 6521 6016 6841 7040
rect 6521 5952 6529 6016
rect 6593 5952 6609 6016
rect 6673 5952 6689 6016
rect 6753 5952 6769 6016
rect 6833 5952 6841 6016
rect 6521 5556 6841 5952
rect 6521 5320 6563 5556
rect 6799 5320 6841 5556
rect 6521 4928 6841 5320
rect 6521 4864 6529 4928
rect 6593 4864 6609 4928
rect 6673 4864 6689 4928
rect 6753 4864 6769 4928
rect 6833 4864 6841 4928
rect 6521 3840 6841 4864
rect 6521 3776 6529 3840
rect 6593 3776 6609 3840
rect 6673 3776 6689 3840
rect 6753 3776 6769 3840
rect 6833 3776 6841 3840
rect 6521 3381 6841 3776
rect 6521 3145 6563 3381
rect 6799 3145 6841 3381
rect 6521 2752 6841 3145
rect 6521 2688 6529 2752
rect 6593 2688 6609 2752
rect 6673 2688 6689 2752
rect 6753 2688 6769 2752
rect 6833 2688 6841 2752
rect 6521 2128 6841 2688
rect 7181 10912 7501 10928
rect 7181 10848 7189 10912
rect 7253 10848 7269 10912
rect 7333 10848 7349 10912
rect 7413 10848 7429 10912
rect 7493 10848 7501 10912
rect 7181 10566 7501 10848
rect 7181 10330 7223 10566
rect 7459 10330 7501 10566
rect 7181 9824 7501 10330
rect 7181 9760 7189 9824
rect 7253 9760 7269 9824
rect 7333 9760 7349 9824
rect 7413 9760 7429 9824
rect 7493 9760 7501 9824
rect 7181 8736 7501 9760
rect 7181 8672 7189 8736
rect 7253 8672 7269 8736
rect 7333 8672 7349 8736
rect 7413 8672 7429 8736
rect 7493 8672 7501 8736
rect 7181 8391 7501 8672
rect 7181 8155 7223 8391
rect 7459 8155 7501 8391
rect 7181 7648 7501 8155
rect 7181 7584 7189 7648
rect 7253 7584 7269 7648
rect 7333 7584 7349 7648
rect 7413 7584 7429 7648
rect 7493 7584 7501 7648
rect 7181 6560 7501 7584
rect 7181 6496 7189 6560
rect 7253 6496 7269 6560
rect 7333 6496 7349 6560
rect 7413 6496 7429 6560
rect 7493 6496 7501 6560
rect 7181 6216 7501 6496
rect 7181 5980 7223 6216
rect 7459 5980 7501 6216
rect 7181 5472 7501 5980
rect 7181 5408 7189 5472
rect 7253 5408 7269 5472
rect 7333 5408 7349 5472
rect 7413 5408 7429 5472
rect 7493 5408 7501 5472
rect 7181 4384 7501 5408
rect 7181 4320 7189 4384
rect 7253 4320 7269 4384
rect 7333 4320 7349 4384
rect 7413 4320 7429 4384
rect 7493 4320 7501 4384
rect 7181 4041 7501 4320
rect 7181 3805 7223 4041
rect 7459 3805 7501 4041
rect 7181 3296 7501 3805
rect 7181 3232 7189 3296
rect 7253 3232 7269 3296
rect 7333 3232 7349 3296
rect 7413 3232 7429 3296
rect 7493 3232 7501 3296
rect 7181 2208 7501 3232
rect 7181 2144 7189 2208
rect 7253 2144 7269 2208
rect 7333 2144 7349 2208
rect 7413 2144 7429 2208
rect 7493 2144 7501 2208
rect 7181 2128 7501 2144
rect 8752 10368 9072 10928
rect 8752 10304 8760 10368
rect 8824 10304 8840 10368
rect 8904 10304 8920 10368
rect 8984 10304 9000 10368
rect 9064 10304 9072 10368
rect 8752 9906 9072 10304
rect 8752 9670 8794 9906
rect 9030 9670 9072 9906
rect 8752 9280 9072 9670
rect 8752 9216 8760 9280
rect 8824 9216 8840 9280
rect 8904 9216 8920 9280
rect 8984 9216 9000 9280
rect 9064 9216 9072 9280
rect 8752 8192 9072 9216
rect 8752 8128 8760 8192
rect 8824 8128 8840 8192
rect 8904 8128 8920 8192
rect 8984 8128 9000 8192
rect 9064 8128 9072 8192
rect 8752 7731 9072 8128
rect 8752 7495 8794 7731
rect 9030 7495 9072 7731
rect 8752 7104 9072 7495
rect 8752 7040 8760 7104
rect 8824 7040 8840 7104
rect 8904 7040 8920 7104
rect 8984 7040 9000 7104
rect 9064 7040 9072 7104
rect 8752 6016 9072 7040
rect 8752 5952 8760 6016
rect 8824 5952 8840 6016
rect 8904 5952 8920 6016
rect 8984 5952 9000 6016
rect 9064 5952 9072 6016
rect 8752 5556 9072 5952
rect 8752 5320 8794 5556
rect 9030 5320 9072 5556
rect 8752 4928 9072 5320
rect 8752 4864 8760 4928
rect 8824 4864 8840 4928
rect 8904 4864 8920 4928
rect 8984 4864 9000 4928
rect 9064 4864 9072 4928
rect 8752 3840 9072 4864
rect 8752 3776 8760 3840
rect 8824 3776 8840 3840
rect 8904 3776 8920 3840
rect 8984 3776 9000 3840
rect 9064 3776 9072 3840
rect 8752 3381 9072 3776
rect 8752 3145 8794 3381
rect 9030 3145 9072 3381
rect 8752 2752 9072 3145
rect 8752 2688 8760 2752
rect 8824 2688 8840 2752
rect 8904 2688 8920 2752
rect 8984 2688 9000 2752
rect 9064 2688 9072 2752
rect 8752 2128 9072 2688
rect 9412 10912 9732 10928
rect 9412 10848 9420 10912
rect 9484 10848 9500 10912
rect 9564 10848 9580 10912
rect 9644 10848 9660 10912
rect 9724 10848 9732 10912
rect 9412 10566 9732 10848
rect 9412 10330 9454 10566
rect 9690 10330 9732 10566
rect 9412 9824 9732 10330
rect 9412 9760 9420 9824
rect 9484 9760 9500 9824
rect 9564 9760 9580 9824
rect 9644 9760 9660 9824
rect 9724 9760 9732 9824
rect 9412 8736 9732 9760
rect 9412 8672 9420 8736
rect 9484 8672 9500 8736
rect 9564 8672 9580 8736
rect 9644 8672 9660 8736
rect 9724 8672 9732 8736
rect 9412 8391 9732 8672
rect 9412 8155 9454 8391
rect 9690 8155 9732 8391
rect 9412 7648 9732 8155
rect 9412 7584 9420 7648
rect 9484 7584 9500 7648
rect 9564 7584 9580 7648
rect 9644 7584 9660 7648
rect 9724 7584 9732 7648
rect 9412 6560 9732 7584
rect 9412 6496 9420 6560
rect 9484 6496 9500 6560
rect 9564 6496 9580 6560
rect 9644 6496 9660 6560
rect 9724 6496 9732 6560
rect 9412 6216 9732 6496
rect 9412 5980 9454 6216
rect 9690 5980 9732 6216
rect 9412 5472 9732 5980
rect 9412 5408 9420 5472
rect 9484 5408 9500 5472
rect 9564 5408 9580 5472
rect 9644 5408 9660 5472
rect 9724 5408 9732 5472
rect 9412 4384 9732 5408
rect 9412 4320 9420 4384
rect 9484 4320 9500 4384
rect 9564 4320 9580 4384
rect 9644 4320 9660 4384
rect 9724 4320 9732 4384
rect 9412 4041 9732 4320
rect 9412 3805 9454 4041
rect 9690 3805 9732 4041
rect 9412 3296 9732 3805
rect 9412 3232 9420 3296
rect 9484 3232 9500 3296
rect 9564 3232 9580 3296
rect 9644 3232 9660 3296
rect 9724 3232 9732 3296
rect 9412 2208 9732 3232
rect 9412 2144 9420 2208
rect 9484 2144 9500 2208
rect 9564 2144 9580 2208
rect 9644 2144 9660 2208
rect 9724 2144 9732 2208
rect 9412 2128 9732 2144
<< via4 >>
rect 2101 9670 2337 9906
rect 2101 7495 2337 7731
rect 2101 5320 2337 5556
rect 2101 3145 2337 3381
rect 2761 10330 2997 10566
rect 2761 8155 2997 8391
rect 2761 5980 2997 6216
rect 4332 9670 4568 9906
rect 4332 7495 4568 7731
rect 2761 3805 2997 4041
rect 4332 5320 4568 5556
rect 4332 3145 4568 3381
rect 4992 10330 5228 10566
rect 4992 8155 5228 8391
rect 4992 5980 5228 6216
rect 4992 3805 5228 4041
rect 6563 9670 6799 9906
rect 6563 7495 6799 7731
rect 6563 5320 6799 5556
rect 6563 3145 6799 3381
rect 7223 10330 7459 10566
rect 7223 8155 7459 8391
rect 7223 5980 7459 6216
rect 7223 3805 7459 4041
rect 8794 9670 9030 9906
rect 8794 7495 9030 7731
rect 8794 5320 9030 5556
rect 8794 3145 9030 3381
rect 9454 10330 9690 10566
rect 9454 8155 9690 8391
rect 9454 5980 9690 6216
rect 9454 3805 9690 4041
<< metal5 >>
rect 1056 10566 10076 10608
rect 1056 10330 2761 10566
rect 2997 10330 4992 10566
rect 5228 10330 7223 10566
rect 7459 10330 9454 10566
rect 9690 10330 10076 10566
rect 1056 10288 10076 10330
rect 1056 9906 10076 9948
rect 1056 9670 2101 9906
rect 2337 9670 4332 9906
rect 4568 9670 6563 9906
rect 6799 9670 8794 9906
rect 9030 9670 10076 9906
rect 1056 9628 10076 9670
rect 1056 8391 10076 8433
rect 1056 8155 2761 8391
rect 2997 8155 4992 8391
rect 5228 8155 7223 8391
rect 7459 8155 9454 8391
rect 9690 8155 10076 8391
rect 1056 8113 10076 8155
rect 1056 7731 10076 7773
rect 1056 7495 2101 7731
rect 2337 7495 4332 7731
rect 4568 7495 6563 7731
rect 6799 7495 8794 7731
rect 9030 7495 10076 7731
rect 1056 7453 10076 7495
rect 1056 6216 10076 6258
rect 1056 5980 2761 6216
rect 2997 5980 4992 6216
rect 5228 5980 7223 6216
rect 7459 5980 9454 6216
rect 9690 5980 10076 6216
rect 1056 5938 10076 5980
rect 1056 5556 10076 5598
rect 1056 5320 2101 5556
rect 2337 5320 4332 5556
rect 4568 5320 6563 5556
rect 6799 5320 8794 5556
rect 9030 5320 10076 5556
rect 1056 5278 10076 5320
rect 1056 4041 10076 4083
rect 1056 3805 2761 4041
rect 2997 3805 4992 4041
rect 5228 3805 7223 4041
rect 7459 3805 9454 4041
rect 9690 3805 10076 4041
rect 1056 3763 10076 3805
rect 1056 3381 10076 3423
rect 1056 3145 2101 3381
rect 2337 3145 4332 3381
rect 4568 3145 6563 3381
rect 6799 3145 8794 3381
rect 9030 3145 10076 3381
rect 1056 3103 10076 3145
use sky130_fd_sc_hd__inv_2  _072_
timestamp 0
transform -1 0 3496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 0
transform -1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _074_
timestamp 0
transform -1 0 2668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _075_
timestamp 0
transform -1 0 4232 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 0
transform 1 0 4600 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _077_
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 0
transform -1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _079_
timestamp 0
transform 1 0 3864 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 0
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _082_
timestamp 0
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _083_
timestamp 0
transform 1 0 2668 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _084_
timestamp 0
transform -1 0 2668 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _085_
timestamp 0
transform 1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _086_
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 0
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 0
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 0
transform -1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 0
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 0
transform -1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 0
transform 1 0 2208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 0
transform -1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _099_
timestamp 0
transform -1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _100_
timestamp 0
transform 1 0 7452 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _101_
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _102_
timestamp 0
transform 1 0 4784 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _103_
timestamp 0
transform -1 0 5152 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _104_
timestamp 0
transform 1 0 5152 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _105_
timestamp 0
transform -1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _106_
timestamp 0
transform -1 0 7084 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _107_
timestamp 0
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _108_
timestamp 0
transform 1 0 5520 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _109_
timestamp 0
transform -1 0 8004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _110_
timestamp 0
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _111_
timestamp 0
transform 1 0 7452 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _112_
timestamp 0
transform 1 0 6992 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _113_
timestamp 0
transform -1 0 7912 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _114_
timestamp 0
transform -1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _115_
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _116_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _117_
timestamp 0
transform 1 0 4416 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _118_
timestamp 0
transform 1 0 4048 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _119_
timestamp 0
transform -1 0 4784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _120_
timestamp 0
transform 1 0 4140 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _121_
timestamp 0
transform 1 0 4968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _122_
timestamp 0
transform -1 0 5428 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _123_
timestamp 0
transform 1 0 4968 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _124_
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _125_
timestamp 0
transform -1 0 7544 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _126_
timestamp 0
transform -1 0 7360 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _127_
timestamp 0
transform -1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 0
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _129_
timestamp 0
transform -1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _130_
timestamp 0
transform -1 0 6992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _131_
timestamp 0
transform -1 0 7360 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _132_
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _133_
timestamp 0
transform 1 0 4968 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 0
transform -1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _135_
timestamp 0
transform 1 0 7268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 0
transform -1 0 8096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _137_
timestamp 0
transform -1 0 2484 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 0
transform -1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _139_
timestamp 0
transform 1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 0
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 0
transform -1 0 5520 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 0
transform -1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _143_
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 0
transform -1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _145_
timestamp 0
transform 1 0 3220 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 0
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _147_
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 0
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _149_
timestamp 0
transform 1 0 2668 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _150_
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _151_
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _152_
timestamp 0
transform 1 0 1564 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _153_
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _154_
timestamp 0
transform 1 0 1472 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _155_
timestamp 0
transform 1 0 1656 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _156_
timestamp 0
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _157_
timestamp 0
transform 1 0 8096 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _158_
timestamp 0
transform 1 0 8280 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _159_
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _160_
timestamp 0
transform 1 0 7268 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _161_
timestamp 0
transform 1 0 5428 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _162_
timestamp 0
transform 1 0 7912 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _163_
timestamp 0
transform 1 0 2116 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _164_
timestamp 0
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _165_
timestamp 0
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _166_
timestamp 0
transform -1 0 5888 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _167_
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _168_
timestamp 0
transform 1 0 8280 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 0
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 0
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 0
transform -1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 0
transform -1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_20
timestamp 0
transform 1 0 2944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_66
timestamp 0
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79
timestamp 0
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_91
timestamp 0
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 0
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_83
timestamp 0
transform 1 0 8740 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_90
timestamp 0
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_9
timestamp 0
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_40
timestamp 0
transform 1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_73
timestamp 0
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 0
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_18
timestamp 0
transform 1 0 2760 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_40
timestamp 0
transform 1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_68
timestamp 0
transform 1 0 7360 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_76
timestamp 0
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 0
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_40
timestamp 0
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_59
timestamp 0
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_63
timestamp 0
transform 1 0 6900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_74
timestamp 0
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_17
timestamp 0
transform 1 0 2668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_29
timestamp 0
transform 1 0 3772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_36
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_37
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_49
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_72
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 0
transform 1 0 8096 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_93
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_28
timestamp 0
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_66
timestamp 0
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_74
timestamp 0
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_92
timestamp 0
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_23
timestamp 0
transform 1 0 3220 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 0
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_68
timestamp 0
transform 1 0 7360 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_48
timestamp 0
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_12
timestamp 0
transform 1 0 2208 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_43
timestamp 0
transform 1 0 5060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_51
timestamp 0
transform 1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_57
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_68
timestamp 0
transform 1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 0
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_10
timestamp 0
transform 1 0 2024 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_49
timestamp 0
transform 1 0 5612 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_23
timestamp 0
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_28
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_36
timestamp 0
transform 1 0 4416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_48
timestamp 0
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 0
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_70
timestamp 0
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_26
timestamp 0
transform 1 0 3496 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_29
timestamp 0
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_37
timestamp 0
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_63
timestamp 0
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_72
timestamp 0
transform 1 0 7728 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_82
timestamp 0
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_91
timestamp 0
transform 1 0 9476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 3220 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 6256 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 9752 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 4784 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 8832 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform -1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output2
timestamp 0
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output3
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 0
transform -1 0 1932 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 0
transform 1 0 9200 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 0
transform -1 0 7728 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 0
transform -1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 0
transform -1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 0
transform 1 0 8924 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output10
timestamp 0
transform -1 0 9660 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 0
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform 1 0 7268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 0
transform 1 0 9200 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 0
transform -1 0 3680 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform -1 0 3220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 0
transform 1 0 8280 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 0
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 0
transform -1 0 2576 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 0
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 0
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 0
transform -1 0 5336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 0
transform -1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output25
timestamp 0
transform -1 0 8280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 0
transform 1 0 3956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 0
transform -1 0 6900 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output28
timestamp 0
transform 1 0 7820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 0
transform -1 0 1932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 0
transform -1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 10028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 10028 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 10028 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 0
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 0
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5566 10880 5566 10880 4 gnd
rlabel metal1 s 5566 10336 5566 10336 4 vdd
rlabel metal1 s 8694 8840 8694 8840 4 R0[0]
rlabel metal2 s 5842 1520 5842 1520 4 R0[1]
rlabel metal3 s 1096 9588 1096 9588 4 R0[2]
rlabel metal1 s 9798 7718 9798 7718 4 R0[3]
rlabel metal1 s 7222 10778 7222 10778 4 R1[0]
rlabel metal2 s 9062 1520 9062 1520 4 R1[1]
rlabel metal3 s 843 1428 843 1428 4 R1[2]
rlabel metal2 s 9338 11543 9338 11543 4 R1[3]
rlabel metal2 s 9246 9571 9246 9571 4 R2[0]
rlabel metal1 s 9338 4522 9338 4522 4 R2[1]
rlabel metal2 s 46 1792 46 1792 4 R2[2]
rlabel metal2 s 10994 1622 10994 1622 4 R2[3]
rlabel metal1 s 9982 10234 9982 10234 4 R3[0]
rlabel metal2 s 2622 1571 2622 1571 4 R3[1]
rlabel metal2 s 2622 11672 2622 11672 4 R3[2]
rlabel metal3 s 843 4828 843 4828 4 R3[3]
rlabel metal1 s 2622 8432 2622 8432 4 _000_
rlabel metal1 s 6164 8058 6164 8058 4 _001_
rlabel metal1 s 1886 6358 1886 6358 4 _002_
rlabel metal1 s 1932 8398 1932 8398 4 _003_
rlabel metal1 s 3956 8058 3956 8058 4 _004_
rlabel metal1 s 7551 8874 7551 8874 4 _005_
rlabel metal1 s 2997 6358 2997 6358 4 _006_
rlabel metal1 s 3319 8874 3319 8874 4 _007_
rlabel metal1 s 8781 9622 8781 9622 4 _008_
rlabel metal1 s 2157 2414 2157 2414 4 _009_
rlabel metal2 s 2254 9826 2254 9826 4 _010_
rlabel metal2 s 1978 4216 1978 4216 4 _011_
rlabel metal1 s 8316 6290 8316 6290 4 _012_
rlabel metal1 s 8500 4114 8500 4114 4 _013_
rlabel metal1 s 5734 3434 5734 3434 4 _014_
rlabel metal2 s 7585 3026 7585 3026 4 _015_
rlabel metal2 s 5842 9826 5842 9826 4 _016_
rlabel metal1 s 8126 5270 8126 5270 4 _017_
rlabel metal1 s 2060 3502 2060 3502 4 _018_
rlabel metal2 s 7958 9554 7958 9554 4 _019_
rlabel metal1 s 5060 8058 5060 8058 4 _020_
rlabel metal2 s 5570 3026 5570 3026 4 _021_
rlabel metal1 s 3460 5678 3460 5678 4 _022_
rlabel metal1 s 8494 7446 8494 7446 4 _023_
rlabel metal1 s 5152 3502 5152 3502 4 _024_
rlabel metal1 s 4922 3502 4922 3502 4 _025_
rlabel metal1 s 6486 4114 6486 4114 4 _026_
rlabel metal1 s 7268 7854 7268 7854 4 _027_
rlabel metal1 s 6716 6766 6716 6766 4 _028_
rlabel metal1 s 6670 6426 6670 6426 4 _029_
rlabel metal1 s 7084 6834 7084 6834 4 _030_
rlabel metal2 s 7130 4267 7130 4267 4 _031_
rlabel metal1 s 6896 3162 6896 3162 4 _032_
rlabel metal1 s 7406 3536 7406 3536 4 _033_
rlabel metal1 s 5612 9554 5612 9554 4 _034_
rlabel metal1 s 7774 5678 7774 5678 4 _035_
rlabel metal1 s 1518 4080 1518 4080 4 _036_
rlabel metal1 s 8096 8942 8096 8942 4 _037_
rlabel metal1 s 4968 7514 4968 7514 4 _038_
rlabel metal1 s 5382 2448 5382 2448 4 _039_
rlabel metal1 s 4462 6289 4462 6289 4 _040_
rlabel metal1 s 8004 6426 8004 6426 4 _041_
rlabel metal1 s 7636 6290 7636 6290 4 _042_
rlabel metal1 s 6026 5712 6026 5712 4 _043_
rlabel metal1 s 4324 5338 4324 5338 4 _044_
rlabel metal1 s 6118 7922 6118 7922 4 _045_
rlabel metal1 s 2162 6767 2162 6767 4 _046_
rlabel metal1 s 1840 6766 1840 6766 4 _047_
rlabel metal1 s 9108 8330 9108 8330 4 _048_
rlabel metal2 s 3818 3876 3818 3876 4 _049_
rlabel metal2 s 3266 9996 3266 9996 4 _050_
rlabel metal1 s 1794 4182 1794 4182 4 _051_
rlabel metal1 s 8694 6970 8694 6970 4 _052_
rlabel metal2 s 8050 7174 8050 7174 4 _053_
rlabel metal1 s 5244 5882 5244 5882 4 _054_
rlabel metal2 s 4554 6528 4554 6528 4 _055_
rlabel metal2 s 5750 5644 5750 5644 4 _056_
rlabel metal1 s 6348 5338 6348 5338 4 _057_
rlabel metal1 s 6440 5678 6440 5678 4 _058_
rlabel metal2 s 5658 5338 5658 5338 4 _059_
rlabel metal1 s 7038 5168 7038 5168 4 _060_
rlabel metal1 s 7176 5202 7176 5202 4 _061_
rlabel metal1 s 7360 5066 7360 5066 4 _062_
rlabel metal1 s 7774 4794 7774 4794 4 _063_
rlabel metal2 s 7406 4896 7406 4896 4 _064_
rlabel metal2 s 5198 4828 5198 4828 4 _065_
rlabel metal1 s 3910 7310 3910 7310 4 _066_
rlabel metal1 s 4554 7378 4554 7378 4 _067_
rlabel metal1 s 4784 4590 4784 4590 4 _068_
rlabel metal2 s 4738 4522 4738 4522 4 _069_
rlabel metal1 s 4508 4046 4508 4046 4 _070_
rlabel metal1 s 4968 4114 4968 4114 4 _071_
rlabel metal3 s 1303 2788 1303 2788 4 clk
rlabel metal1 s 4508 7446 4508 7446 4 clknet_0_clk
rlabel metal1 s 2162 3638 2162 3638 4 clknet_1_0__leaf_clk
rlabel metal1 s 2714 8534 2714 8534 4 clknet_1_1__leaf_clk
rlabel metal3 s 9622 748 9622 748 4 halt
rlabel metal3 s 820 8228 820 8228 4 instr[0]
rlabel metal2 s 1334 1860 1334 1860 4 instr[1]
rlabel metal2 s 1334 11400 1334 11400 4 instr[2]
rlabel metal1 s 9522 2822 9522 2822 4 instr[3]
rlabel metal2 s 4554 1554 4554 1554 4 instr[4]
rlabel metal3 s 1142 11628 1142 11628 4 instr[5]
rlabel metal1 s 8142 9350 8142 9350 4 instr[6]
rlabel metal1 s 4048 10778 4048 10778 4 instr[7]
rlabel metal1 s 7866 8874 7866 8874 4 net1
rlabel metal1 s 9430 6426 9430 6426 4 net10
rlabel metal1 s 8418 4488 8418 4488 4 net11
rlabel metal1 s 4572 3502 4572 3502 4 net12
rlabel metal1 s 7406 2312 7406 2312 4 net13
rlabel metal1 s 9752 9418 9752 9418 4 net14
rlabel metal1 s 3542 2312 3542 2312 4 net15
rlabel metal1 s 3082 10132 3082 10132 4 net16
rlabel metal1 s 1564 5134 1564 5134 4 net17
rlabel metal2 s 2714 6833 2714 6833 4 net18
rlabel metal1 s 1932 7854 1932 7854 4 net19
rlabel metal1 s 7406 7412 7406 7412 4 net2
rlabel metal1 s 2438 2992 2438 2992 4 net20
rlabel metal1 s 2438 9928 2438 9928 4 net21
rlabel metal1 s 7682 5202 7682 5202 4 net22
rlabel metal1 s 1794 9690 1794 9690 4 net23
rlabel metal1 s 1978 9486 1978 9486 4 net24
rlabel metal1 s 8188 9146 8188 9146 4 net25
rlabel metal1 s 3864 9690 3864 9690 4 net26
rlabel metal1 s 2622 6664 2622 6664 4 net27
rlabel metal1 s 7590 2414 7590 2414 4 net28
rlabel metal1 s 2476 6630 2476 6630 4 net29
rlabel metal1 s 5612 2346 5612 2346 4 net3
rlabel metal2 s 3082 9741 3082 9741 4 net30
rlabel metal1 s 4692 9894 4692 9894 4 net31
rlabel metal1 s 1702 8466 1702 8466 4 net32
rlabel metal2 s 5290 3706 5290 3706 4 net33
rlabel metal1 s 2484 5202 2484 5202 4 net34
rlabel metal1 s 3634 10234 3634 10234 4 net35
rlabel metal1 s 8970 8466 8970 8466 4 net36
rlabel metal1 s 8372 3502 8372 3502 4 net37
rlabel metal1 s 4324 2618 4324 2618 4 net38
rlabel metal1 s 2898 6732 2898 6732 4 net39
rlabel metal2 s 2622 9214 2622 9214 4 net4
rlabel metal1 s 3450 7888 3450 7888 4 net40
rlabel metal1 s 2300 4182 2300 4182 4 net41
rlabel metal2 s 7038 10234 7038 10234 4 net42
rlabel metal1 s 6026 9622 6026 9622 4 net43
rlabel metal1 s 8142 5746 8142 5746 4 net44
rlabel metal1 s 7038 4726 7038 4726 4 net45
rlabel metal1 s 8142 6664 8142 6664 4 net46
rlabel metal1 s 9706 7786 9706 7786 4 net5
rlabel metal1 s 7360 9486 7360 9486 4 net6
rlabel metal1 s 9522 5780 9522 5780 4 net7
rlabel metal1 s 2277 3434 2277 3434 4 net8
rlabel metal1 s 8602 9894 8602 9894 4 net9
rlabel metal1 s 6164 10778 6164 10778 4 pc[0]
rlabel metal2 s 7774 1520 7774 1520 4 pc[1]
rlabel metal3 s 820 6188 820 6188 4 pc[2]
rlabel metal1 s 2254 10744 2254 10744 4 pc[3]
rlabel metal1 s 9844 5270 9844 5270 4 reset
flabel metal3 s 10390 8848 11190 8968 0 FreeSans 600 0 0 0 R0[0]
port 1 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 R0[1]
port 2 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 R0[2]
port 3 nsew
flabel metal3 s 10390 7488 11190 7608 0 FreeSans 600 0 0 0 R0[3]
port 4 nsew
flabel metal2 s 7102 12534 7158 13334 0 FreeSans 280 90 0 0 R1[0]
port 5 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 R1[1]
port 6 nsew
flabel metal3 s 0 1368 800 1488 0 FreeSans 600 0 0 0 R1[2]
port 7 nsew
flabel metal3 s 10390 12248 11190 12368 0 FreeSans 600 0 0 0 R1[3]
port 8 nsew
flabel metal2 s 9034 12534 9090 13334 0 FreeSans 280 90 0 0 R2[0]
port 9 nsew
flabel metal3 s 10390 4088 11190 4208 0 FreeSans 600 0 0 0 R2[1]
port 10 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 R2[2]
port 11 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 R2[3]
port 12 nsew
flabel metal2 s 10322 12534 10378 13334 0 FreeSans 280 90 0 0 R3[0]
port 13 nsew
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 R3[1]
port 14 nsew
flabel metal2 s 2594 12534 2650 13334 0 FreeSans 280 90 0 0 R3[2]
port 15 nsew
flabel metal3 s 0 4768 800 4888 0 FreeSans 600 0 0 0 R3[3]
port 16 nsew
flabel metal3 s 0 2728 800 2848 0 FreeSans 600 0 0 0 clk
port 17 nsew
flabel metal5 s 1056 10288 10076 10608 0 FreeSans 3200 0 0 0 gnd
port 18 nsew
flabel metal5 s 1056 8113 10076 8433 0 FreeSans 3200 0 0 0 gnd
port 18 nsew
flabel metal5 s 1056 5938 10076 6258 0 FreeSans 3200 0 0 0 gnd
port 18 nsew
flabel metal5 s 1056 3763 10076 4083 0 FreeSans 3200 0 0 0 gnd
port 18 nsew
flabel metal4 s 9412 2128 9732 10928 0 FreeSans 2400 90 0 0 gnd
port 18 nsew
flabel metal4 s 7181 2128 7501 10928 0 FreeSans 2400 90 0 0 gnd
port 18 nsew
flabel metal4 s 4950 2128 5270 10928 0 FreeSans 2400 90 0 0 gnd
port 18 nsew
flabel metal4 s 2719 2128 3039 10928 0 FreeSans 2400 90 0 0 gnd
port 18 nsew
flabel metal3 s 10390 688 11190 808 0 FreeSans 600 0 0 0 halt
port 19 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 instr[0]
port 20 nsew
flabel metal2 s 1306 0 1362 800 0 FreeSans 280 90 0 0 instr[1]
port 21 nsew
flabel metal2 s 1306 12534 1362 13334 0 FreeSans 280 90 0 0 instr[2]
port 22 nsew
flabel metal3 s 10390 2728 11190 2848 0 FreeSans 600 0 0 0 instr[3]
port 23 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 instr[4]
port 24 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 instr[5]
port 25 nsew
flabel metal3 s 10390 10888 11190 11008 0 FreeSans 600 0 0 0 instr[6]
port 26 nsew
flabel metal2 s 3882 12534 3938 13334 0 FreeSans 280 90 0 0 instr[7]
port 27 nsew
flabel metal2 s 5814 12534 5870 13334 0 FreeSans 280 90 0 0 pc[0]
port 28 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 pc[1]
port 29 nsew
flabel metal3 s 0 6128 800 6248 0 FreeSans 600 0 0 0 pc[2]
port 30 nsew
flabel metal3 s 0 12928 800 13048 0 FreeSans 600 0 0 0 pc[3]
port 31 nsew
flabel metal3 s 10390 5448 11190 5568 0 FreeSans 600 0 0 0 reset
port 32 nsew
flabel metal5 s 1056 9628 10076 9948 0 FreeSans 3200 0 0 0 vdd
port 33 nsew
flabel metal5 s 1056 7453 10076 7773 0 FreeSans 3200 0 0 0 vdd
port 33 nsew
flabel metal5 s 1056 5278 10076 5598 0 FreeSans 3200 0 0 0 vdd
port 33 nsew
flabel metal5 s 1056 3103 10076 3423 0 FreeSans 3200 0 0 0 vdd
port 33 nsew
flabel metal4 s 8752 2128 9072 10928 0 FreeSans 2400 90 0 0 vdd
port 33 nsew
flabel metal4 s 6521 2128 6841 10928 0 FreeSans 2400 90 0 0 vdd
port 33 nsew
flabel metal4 s 4290 2128 4610 10928 0 FreeSans 2400 90 0 0 vdd
port 33 nsew
flabel metal4 s 2059 2128 2379 10928 0 FreeSans 2400 90 0 0 vdd
port 33 nsew
<< properties >>
string FIXED_BBOX 0 0 11190 13334
<< end >>
