VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO riscv32
  CLASS BLOCK ;
  FOREIGN riscv32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 55.950 BY 66.670 ;
  PIN R0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 51.950 44.240 55.950 44.840 ;
    END
  END R0[0]
  PIN R0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END R0[1]
  PIN R0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END R0[2]
  PIN R0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 37.440 55.950 38.040 ;
    END
  END R0[3]
  PIN R1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 62.670 35.790 66.670 ;
    END
  END R1[0]
  PIN R1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END R1[1]
  PIN R1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END R1[2]
  PIN R1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 61.240 55.950 61.840 ;
    END
  END R1[3]
  PIN R2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 62.670 45.450 66.670 ;
    END
  END R2[0]
  PIN R2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 20.440 55.950 21.040 ;
    END
  END R2[1]
  PIN R2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END R2[2]
  PIN R2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END R2[3]
  PIN R3[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 62.670 51.890 66.670 ;
    END
  END R3[0]
  PIN R3[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END R3[1]
  PIN R3[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.970 62.670 13.250 66.670 ;
    END
  END R3[2]
  PIN R3[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END R3[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END clk
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.595 10.640 15.195 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.750 10.640 26.350 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.905 10.640 37.505 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.060 10.640 48.660 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.815 50.380 20.415 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.690 50.380 31.290 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.565 50.380 42.165 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 51.440 50.380 53.040 ;
    END
  END gnd
  PIN halt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 3.440 55.950 4.040 ;
    END
  END halt
  PIN instr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END instr[0]
  PIN instr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END instr[1]
  PIN instr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 62.670 6.810 66.670 ;
    END
  END instr[2]
  PIN instr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 13.640 55.950 14.240 ;
    END
  END instr[3]
  PIN instr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END instr[4]
  PIN instr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END instr[5]
  PIN instr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 51.950 54.440 55.950 55.040 ;
    END
  END instr[6]
  PIN instr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 62.670 19.690 66.670 ;
    END
  END instr[7]
  PIN pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 29.070 62.670 29.350 66.670 ;
    END
  END pc[0]
  PIN pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END pc[1]
  PIN pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END pc[2]
  PIN pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END pc[3]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 51.950 27.240 55.950 27.840 ;
    END
  END reset
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.295 10.640 11.895 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.450 10.640 23.050 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.605 10.640 34.205 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.760 10.640 45.360 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.515 50.380 17.115 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.390 50.380 27.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.265 50.380 38.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 48.140 50.380 49.740 ;
    END
  END vdd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 50.140 54.485 ;
      LAYER met1 ;
        RECT 0.070 10.640 55.130 54.640 ;
      LAYER met2 ;
        RECT 0.100 62.390 6.250 65.125 ;
        RECT 7.090 62.390 12.690 65.125 ;
        RECT 13.530 62.390 19.130 65.125 ;
        RECT 19.970 62.390 28.790 65.125 ;
        RECT 29.630 62.390 35.230 65.125 ;
        RECT 36.070 62.390 44.890 65.125 ;
        RECT 45.730 62.390 51.330 65.125 ;
        RECT 52.170 62.390 55.100 65.125 ;
        RECT 0.100 4.280 55.100 62.390 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 54.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 64.240 51.950 65.105 ;
        RECT 4.000 62.240 51.950 64.240 ;
        RECT 4.000 60.840 51.550 62.240 ;
        RECT 4.000 58.840 51.950 60.840 ;
        RECT 4.400 57.440 51.950 58.840 ;
        RECT 4.000 55.440 51.950 57.440 ;
        RECT 4.000 54.040 51.550 55.440 ;
        RECT 4.000 48.640 51.950 54.040 ;
        RECT 4.400 47.240 51.950 48.640 ;
        RECT 4.000 45.240 51.950 47.240 ;
        RECT 4.000 43.840 51.550 45.240 ;
        RECT 4.000 41.840 51.950 43.840 ;
        RECT 4.400 40.440 51.950 41.840 ;
        RECT 4.000 38.440 51.950 40.440 ;
        RECT 4.000 37.040 51.550 38.440 ;
        RECT 4.000 31.640 51.950 37.040 ;
        RECT 4.400 30.240 51.950 31.640 ;
        RECT 4.000 28.240 51.950 30.240 ;
        RECT 4.000 26.840 51.550 28.240 ;
        RECT 4.000 24.840 51.950 26.840 ;
        RECT 4.400 23.440 51.950 24.840 ;
        RECT 4.000 21.440 51.950 23.440 ;
        RECT 4.000 20.040 51.550 21.440 ;
        RECT 4.000 14.640 51.950 20.040 ;
        RECT 4.400 13.240 51.550 14.640 ;
        RECT 4.000 7.840 51.950 13.240 ;
        RECT 4.400 6.440 51.950 7.840 ;
        RECT 4.000 4.440 51.950 6.440 ;
        RECT 4.000 3.575 51.550 4.440 ;
      LAYER met4 ;
        RECT 18.695 14.455 19.025 28.385 ;
  END
END riscv32
END LIBRARY

